module star (
input_R1,output_R1,
/*input_R2,output_R2,
input_R3,output_R3,
input_R4,output_R4,
input_R5,output_R5,
input_R6,output_R6,
input_R7,output_R7,
input_R8,output_R8,
input_R9,output_R9,
input_R10,output_R10,
input_R11,output_R11,
input_R12,output_R12,
input_R13,output_R13,
input_R14,output_R14,
input_R15,output_R15,
input_R16,output_R16,
input_R17,output_R17,
input_R18,output_R18,
input_R19,output_R19,
input_R20,output_R20,
input_R21,output_R21,
input_R22,output_R22,
input_R23,output_R23,
input_R24,output_R24,
input_R25,output_R25,
input_R26,output_R26,
input_R27,output_R27,
input_R28,output_R28,
input_R29,output_R29,
input_R30,output_R30,
input_R31,output_R31,
input_R32,output_R32,
input_R33,output_R33,
input_R34,output_R34,
input_R35,output_R35,
input_R36,output_R36,
input_R37,output_R37,
input_R38,output_R38,
input_R39,output_R39,
input_R40,output_R40,
input_R41,output_R41,
input_R42,output_R42,
input_R43,output_R43,
input_R44,output_R44,
input_R45,output_R45,
input_R46,output_R46,
input_R47,output_R47,
input_R48,output_R48,
input_R49,output_R49,
input_R50,output_R50,
input_R51,output_R51,
input_R52,output_R52,
input_R53,output_R53,
input_R54,output_R54,
input_R55,output_R55,
input_R56,output_R56,
input_R57,output_R57,
input_R58,output_R58,
input_R59,output_R59,
input_R60,output_R60,
input_R61,output_R61,
input_R62,output_R62, */
input_R63,output_R63,
clk, rst,  Write, Read);
input clk, rst, Write, Read; 
parameter DATAWID = 8;
input [DATAWID-1:0] input_R1;
output [DATAWID-1:0] output_R1;
wire [DATAWID-1:0] input_R2;
wire [DATAWID-1:0] output_R2;
wire [DATAWID-1:0] input_R3;
wire [DATAWID-1:0] output_R3;
wire [DATAWID-1:0] input_R4;
wire [DATAWID-1:0] output_R4;
wire [DATAWID-1:0] input_R5;
wire [DATAWID-1:0] output_R5;
wire [DATAWID-1:0] input_R6;
wire [DATAWID-1:0] output_R6;
wire [DATAWID-1:0] input_R7;
wire [DATAWID-1:0] output_R7;
wire [DATAWID-1:0] input_R8;
wire [DATAWID-1:0] output_R8;
wire [DATAWID-1:0] input_R9;
wire [DATAWID-1:0] output_R9;
wire [DATAWID-1:0] input_R10;
wire [DATAWID-1:0] output_R10;
wire [DATAWID-1:0] input_R11;
wire [DATAWID-1:0] output_R11;
wire [DATAWID-1:0] input_R12;
wire [DATAWID-1:0] output_R12;
wire [DATAWID-1:0] input_R13;
wire [DATAWID-1:0] output_R13;
wire [DATAWID-1:0] input_R14;
wire [DATAWID-1:0] output_R14;
wire [DATAWID-1:0] input_R15;
wire [DATAWID-1:0] output_R15;
wire [DATAWID-1:0] input_R16;
wire [DATAWID-1:0] output_R16;
wire [DATAWID-1:0] input_R17;
wire [DATAWID-1:0] output_R17;
wire [DATAWID-1:0] input_R18;
wire [DATAWID-1:0] output_R18;
wire [DATAWID-1:0] input_R19;
wire [DATAWID-1:0] output_R19;
wire [DATAWID-1:0] input_R20;
wire [DATAWID-1:0] output_R20;
wire [DATAWID-1:0] input_R21;
wire [DATAWID-1:0] output_R21;
wire [DATAWID-1:0] input_R22;
wire [DATAWID-1:0] output_R22;
wire [DATAWID-1:0] input_R23;
wire [DATAWID-1:0] output_R23;
wire [DATAWID-1:0] input_R24;
wire [DATAWID-1:0] output_R24;
wire [DATAWID-1:0] input_R25;
wire [DATAWID-1:0] output_R25;
wire [DATAWID-1:0] input_R26;
wire [DATAWID-1:0] output_R26;
wire [DATAWID-1:0] input_R27;
wire [DATAWID-1:0] output_R27;
wire [DATAWID-1:0] input_R28;
wire [DATAWID-1:0] output_R28;
wire [DATAWID-1:0] input_R29;
wire [DATAWID-1:0] output_R29;
wire [DATAWID-1:0] input_R30;
wire [DATAWID-1:0] output_R30;
wire [DATAWID-1:0] input_R31;
wire [DATAWID-1:0] output_R31;
wire [DATAWID-1:0] input_R32;
wire [DATAWID-1:0] output_R32;
wire [DATAWID-1:0] input_R33;
wire [DATAWID-1:0] output_R33;
wire [DATAWID-1:0] input_R34;
wire [DATAWID-1:0] output_R34;
wire [DATAWID-1:0] input_R35;
wire [DATAWID-1:0] output_R35;
wire [DATAWID-1:0] input_R36;
wire [DATAWID-1:0] output_R36;
wire [DATAWID-1:0] input_R37;
wire [DATAWID-1:0] output_R37;
wire [DATAWID-1:0] input_R38;
wire [DATAWID-1:0] output_R38;
wire [DATAWID-1:0] input_R39;
wire [DATAWID-1:0] output_R39;
wire [DATAWID-1:0] input_R40;
wire [DATAWID-1:0] output_R40;
wire [DATAWID-1:0] input_R41;
wire [DATAWID-1:0] output_R41;
wire [DATAWID-1:0] input_R42;
wire [DATAWID-1:0] output_R42;
wire [DATAWID-1:0] input_R43;
wire [DATAWID-1:0] output_R43;
wire [DATAWID-1:0] input_R44;
wire [DATAWID-1:0] output_R44;
wire [DATAWID-1:0] input_R45;
wire [DATAWID-1:0] output_R45;
wire [DATAWID-1:0] input_R46;
wire [DATAWID-1:0] output_R46;
wire [DATAWID-1:0] input_R47;
wire [DATAWID-1:0] output_R47;
wire [DATAWID-1:0] input_R48;
wire [DATAWID-1:0] output_R48;
wire [DATAWID-1:0] input_R49;
wire [DATAWID-1:0] output_R49;
wire [DATAWID-1:0] input_R50;
wire [DATAWID-1:0] output_R50;
wire [DATAWID-1:0] input_R51;
wire [DATAWID-1:0] output_R51;
wire [DATAWID-1:0] input_R52;
wire [DATAWID-1:0] output_R52;
wire [DATAWID-1:0] input_R53;
wire [DATAWID-1:0] output_R53;
wire [DATAWID-1:0] input_R54;
wire [DATAWID-1:0] output_R54;
wire [DATAWID-1:0] input_R55;
wire [DATAWID-1:0] output_R55;
wire [DATAWID-1:0] input_R56;
wire [DATAWID-1:0] output_R56;
wire [DATAWID-1:0] input_R57;
wire [DATAWID-1:0] output_R57;
wire [DATAWID-1:0] input_R58;
wire [DATAWID-1:0] output_R58;
wire [DATAWID-1:0] input_R59;
wire [DATAWID-1:0] output_R59;
wire [DATAWID-1:0] input_R60;
wire [DATAWID-1:0] output_R60;
wire [DATAWID-1:0] input_R61;
wire [DATAWID-1:0] output_R61;
wire [DATAWID-1:0] input_R62;
wire [DATAWID-1:0] output_R62;
input [DATAWID-1:0] input_R63;
output [DATAWID-1:0] output_R63;
reg [DATAWID-1:0] R0_in0;
wire [DATAWID-1:0] R0_out0;
reg [DATAWID-1:0] R0_in1;
wire [DATAWID-1:0] R0_out1;
reg [DATAWID-1:0] R0_in2;
wire [DATAWID-1:0] R0_out2;
reg [DATAWID-1:0] R0_in3;
wire [DATAWID-1:0] R0_out3;
reg [DATAWID-1:0] R0_in4;
wire [DATAWID-1:0] R0_out4;
reg [DATAWID-1:0] R0_in5;
wire [DATAWID-1:0] R0_out5;
reg [DATAWID-1:0] R0_in6;
wire [DATAWID-1:0] R0_out6;
reg [DATAWID-1:0] R0_in7;
wire [DATAWID-1:0] R0_out7;
reg [DATAWID-1:0] R0_in8;
wire [DATAWID-1:0] R0_out8;
reg [DATAWID-1:0] R0_in9;
wire [DATAWID-1:0] R0_out9;
reg [DATAWID-1:0] R0_in10;
wire [DATAWID-1:0] R0_out10;
reg [DATAWID-1:0] R0_in11;
wire [DATAWID-1:0] R0_out11;
reg [DATAWID-1:0] R0_in12;
wire [DATAWID-1:0] R0_out12;
reg [DATAWID-1:0] R0_in13;
wire [DATAWID-1:0] R0_out13;
reg [DATAWID-1:0] R0_in14;
wire [DATAWID-1:0] R0_out14;
reg [DATAWID-1:0] R0_in15;
wire [DATAWID-1:0] R0_out15;
reg [DATAWID-1:0] R0_in16;
wire [DATAWID-1:0] R0_out16;
reg [DATAWID-1:0] R0_in17;
wire [DATAWID-1:0] R0_out17;
reg [DATAWID-1:0] R0_in18;
wire [DATAWID-1:0] R0_out18;
reg [DATAWID-1:0] R0_in19;
wire [DATAWID-1:0] R0_out19;
reg [DATAWID-1:0] R0_in20;
wire [DATAWID-1:0] R0_out20;
reg [DATAWID-1:0] R0_in21;
wire [DATAWID-1:0] R0_out21;
reg [DATAWID-1:0] R0_in22;
wire [DATAWID-1:0] R0_out22;
reg [DATAWID-1:0] R0_in23;
wire [DATAWID-1:0] R0_out23;
reg [DATAWID-1:0] R0_in24;
wire [DATAWID-1:0] R0_out24;
reg [DATAWID-1:0] R0_in25;
wire [DATAWID-1:0] R0_out25;
reg [DATAWID-1:0] R0_in26;
wire [DATAWID-1:0] R0_out26;
reg [DATAWID-1:0] R0_in27;
wire [DATAWID-1:0] R0_out27;
reg [DATAWID-1:0] R0_in28;
wire [DATAWID-1:0] R0_out28;
reg [DATAWID-1:0] R0_in29;
wire [DATAWID-1:0] R0_out29;
reg [DATAWID-1:0] R0_in30;
wire [DATAWID-1:0] R0_out30;
reg [DATAWID-1:0] R0_in31;
wire [DATAWID-1:0] R0_out31;
reg [DATAWID-1:0] R0_in32;
wire [DATAWID-1:0] R0_out32;
reg [DATAWID-1:0] R0_in33;
wire [DATAWID-1:0] R0_out33;
reg [DATAWID-1:0] R0_in34;
wire [DATAWID-1:0] R0_out34;
reg [DATAWID-1:0] R0_in35;
wire [DATAWID-1:0] R0_out35;
reg [DATAWID-1:0] R0_in36;
wire [DATAWID-1:0] R0_out36;
reg [DATAWID-1:0] R0_in37;
wire [DATAWID-1:0] R0_out37;
reg [DATAWID-1:0] R0_in38;
wire [DATAWID-1:0] R0_out38;
reg [DATAWID-1:0] R0_in39;
wire [DATAWID-1:0] R0_out39;
reg [DATAWID-1:0] R0_in40;
wire [DATAWID-1:0] R0_out40;
reg [DATAWID-1:0] R0_in41;
wire [DATAWID-1:0] R0_out41;
reg [DATAWID-1:0] R0_in42;
wire [DATAWID-1:0] R0_out42;
reg [DATAWID-1:0] R0_in43;
wire [DATAWID-1:0] R0_out43;
reg [DATAWID-1:0] R0_in44;
wire [DATAWID-1:0] R0_out44;
reg [DATAWID-1:0] R0_in45;
wire [DATAWID-1:0] R0_out45;
reg [DATAWID-1:0] R0_in46;
wire [DATAWID-1:0] R0_out46;
reg [DATAWID-1:0] R0_in47;
wire [DATAWID-1:0] R0_out47;
reg [DATAWID-1:0] R0_in48;
wire [DATAWID-1:0] R0_out48;
reg [DATAWID-1:0] R0_in49;
wire [DATAWID-1:0] R0_out49;
reg [DATAWID-1:0] R0_in50;
wire [DATAWID-1:0] R0_out50;
reg [DATAWID-1:0] R0_in51;
wire [DATAWID-1:0] R0_out51;
reg [DATAWID-1:0] R0_in52;
wire [DATAWID-1:0] R0_out52;
reg [DATAWID-1:0] R0_in53;
wire [DATAWID-1:0] R0_out53;
reg [DATAWID-1:0] R0_in54;
wire [DATAWID-1:0] R0_out54;
reg [DATAWID-1:0] R0_in55;
wire [DATAWID-1:0] R0_out55;
reg [DATAWID-1:0] R0_in56;
wire [DATAWID-1:0] R0_out56;
reg [DATAWID-1:0] R0_in57;
wire [DATAWID-1:0] R0_out57;
reg [DATAWID-1:0] R0_in58;
wire [DATAWID-1:0] R0_out58;
reg [DATAWID-1:0] R0_in59;
wire [DATAWID-1:0] R0_out59;
reg [DATAWID-1:0] R0_in60;
wire [DATAWID-1:0] R0_out60;
reg [DATAWID-1:0] R0_in61;
wire [DATAWID-1:0] R0_out61;
reg [DATAWID-1:0] R0_in62;
wire [DATAWID-1:0] R0_out62;
reg [DATAWID-1:0] port1_inR1;
reg [DATAWID-1:0] port1_inR2;
reg [DATAWID-1:0] port1_inR3;
reg [DATAWID-1:0] port1_inR4;
reg [DATAWID-1:0] port1_inR5;
reg [DATAWID-1:0] port1_inR6;
reg [DATAWID-1:0] port1_inR7;
reg [DATAWID-1:0] port1_inR8;
reg [DATAWID-1:0] port1_inR9;
reg [DATAWID-1:0] port1_inR10;
reg [DATAWID-1:0] port1_inR11;
reg [DATAWID-1:0] port1_inR12;
reg [DATAWID-1:0] port1_inR13;
reg [DATAWID-1:0] port1_inR14;
reg [DATAWID-1:0] port1_inR15;
reg [DATAWID-1:0] port1_inR16;
reg [DATAWID-1:0] port1_inR17;
reg [DATAWID-1:0] port1_inR18;
reg [DATAWID-1:0] port1_inR19;
reg [DATAWID-1:0] port1_inR20;
reg [DATAWID-1:0] port1_inR21;
reg [DATAWID-1:0] port1_inR22;
reg [DATAWID-1:0] port1_inR23;
reg [DATAWID-1:0] port1_inR24;
reg [DATAWID-1:0] port1_inR25;
reg [DATAWID-1:0] port1_inR26;
reg [DATAWID-1:0] port1_inR27;
reg [DATAWID-1:0] port1_inR28;
reg [DATAWID-1:0] port1_inR29;
reg [DATAWID-1:0] port1_inR30;
reg [DATAWID-1:0] port1_inR31;
reg [DATAWID-1:0] port1_inR32;
reg [DATAWID-1:0] port1_inR33;
reg [DATAWID-1:0] port1_inR34;
reg [DATAWID-1:0] port1_inR35;
reg [DATAWID-1:0] port1_inR36;
reg [DATAWID-1:0] port1_inR37;
reg [DATAWID-1:0] port1_inR38;
reg [DATAWID-1:0] port1_inR39;
reg [DATAWID-1:0] port1_inR40;
reg [DATAWID-1:0] port1_inR41;
reg [DATAWID-1:0] port1_inR42;
reg [DATAWID-1:0] port1_inR43;
reg [DATAWID-1:0] port1_inR44;
reg [DATAWID-1:0] port1_inR45;
reg [DATAWID-1:0] port1_inR46;
reg [DATAWID-1:0] port1_inR47;
reg [DATAWID-1:0] port1_inR48;
reg [DATAWID-1:0] port1_inR49;
reg [DATAWID-1:0] port1_inR50;
reg [DATAWID-1:0] port1_inR51;
reg [DATAWID-1:0] port1_inR52;
reg [DATAWID-1:0] port1_inR53;
reg [DATAWID-1:0] port1_inR54;
reg [DATAWID-1:0] port1_inR55;
reg [DATAWID-1:0] port1_inR56;
reg [DATAWID-1:0] port1_inR57;
reg [DATAWID-1:0] port1_inR58;
reg [DATAWID-1:0] port1_inR59;
reg [DATAWID-1:0] port1_inR60;
reg [DATAWID-1:0] port1_inR61;
reg [DATAWID-1:0] port1_inR62;
reg [DATAWID-1:0] port1_inR63;
wire [DATAWID-1:0] port1_outR1;
wire [DATAWID-1:0] port1_outR2;
wire [DATAWID-1:0] port1_outR3;
wire [DATAWID-1:0] port1_outR4;
wire [DATAWID-1:0] port1_outR5;
wire [DATAWID-1:0] port1_outR6;
wire [DATAWID-1:0] port1_outR7;
wire [DATAWID-1:0] port1_outR8;
wire [DATAWID-1:0] port1_outR9;
wire [DATAWID-1:0] port1_outR10;
wire [DATAWID-1:0] port1_outR11;
wire [DATAWID-1:0] port1_outR12;
wire [DATAWID-1:0] port1_outR13;
wire [DATAWID-1:0] port1_outR14;
wire [DATAWID-1:0] port1_outR15;
wire [DATAWID-1:0] port1_outR16;
wire [DATAWID-1:0] port1_outR17;
wire [DATAWID-1:0] port1_outR18;
wire [DATAWID-1:0] port1_outR19;
wire [DATAWID-1:0] port1_outR20;
wire [DATAWID-1:0] port1_outR21;
wire [DATAWID-1:0] port1_outR22;
wire [DATAWID-1:0] port1_outR23;
wire [DATAWID-1:0] port1_outR24;
wire [DATAWID-1:0] port1_outR25;
wire [DATAWID-1:0] port1_outR26;
wire [DATAWID-1:0] port1_outR27;
wire [DATAWID-1:0] port1_outR28;
wire [DATAWID-1:0] port1_outR29;
wire [DATAWID-1:0] port1_outR30;
wire [DATAWID-1:0] port1_outR31;
wire [DATAWID-1:0] port1_outR32;
wire [DATAWID-1:0] port1_outR33;
wire [DATAWID-1:0] port1_outR34;
wire [DATAWID-1:0] port1_outR35;
wire [DATAWID-1:0] port1_outR36;
wire [DATAWID-1:0] port1_outR37;
wire [DATAWID-1:0] port1_outR38;
wire [DATAWID-1:0] port1_outR39;
wire [DATAWID-1:0] port1_outR40;
wire [DATAWID-1:0] port1_outR41;
wire [DATAWID-1:0] port1_outR42;
wire [DATAWID-1:0] port1_outR43;
wire [DATAWID-1:0] port1_outR44;
wire [DATAWID-1:0] port1_outR45;
wire [DATAWID-1:0] port1_outR46;
wire [DATAWID-1:0] port1_outR47;
wire [DATAWID-1:0] port1_outR48;
wire [DATAWID-1:0] port1_outR49;
wire [DATAWID-1:0] port1_outR50;
wire [DATAWID-1:0] port1_outR51;
wire [DATAWID-1:0] port1_outR52;
wire [DATAWID-1:0] port1_outR53;
wire [DATAWID-1:0] port1_outR54;
wire [DATAWID-1:0] port1_outR55;
wire [DATAWID-1:0] port1_outR56;
wire [DATAWID-1:0] port1_outR57;
wire [DATAWID-1:0] port1_outR58;
wire [DATAWID-1:0] port1_outR59;
wire [DATAWID-1:0] port1_outR60;
wire [DATAWID-1:0] port1_outR61;
wire [DATAWID-1:0] port1_outR62;
wire [DATAWID-1:0] port1_outR63;
router0 r
( .clk(clk), .rst(reset),
.i000(R0_in0),
.i010(R0_out0),
.i001(R0_in1),
.i011(R0_out1),
.i002(R0_in2),
.i012(R0_out2),
.i003(R0_in3),
.i013(R0_out3),
.i004(R0_in4),
.i014(R0_out4),
.i005(R0_in5),
.i015(R0_out5),
.i006(R0_in6),
.i016(R0_out6),
.i007(R0_in7),
.i017(R0_out7),
.i008(R0_in8),
.i018(R0_out8),
.i009(R0_in9),
.i019(R0_out9),
.i0010(R0_in10),
.i0110(R0_out10),
.i0011(R0_in11),
.i0111(R0_out11),
.i0012(R0_in12),
.i0112(R0_out12),
.i0013(R0_in13),
.i0113(R0_out13),
.i0014(R0_in14),
.i0114(R0_out14),
.i0015(R0_in15),
.i0115(R0_out15),
.i0016(R0_in16),
.i0116(R0_out16),
.i0017(R0_in17),
.i0117(R0_out17),
.i0018(R0_in18),
.i0118(R0_out18),
.i0019(R0_in19),
.i0119(R0_out19),
.i0020(R0_in20),
.i0120(R0_out20),
.i0021(R0_in21),
.i0121(R0_out21),
.i0022(R0_in22),
.i0122(R0_out22),
.i0023(R0_in23),
.i0123(R0_out23),
.i0024(R0_in24),
.i0124(R0_out24),
.i0025(R0_in25),
.i0125(R0_out25),
.i0026(R0_in26),
.i0126(R0_out26),
.i0027(R0_in27),
.i0127(R0_out27),
.i0028(R0_in28),
.i0128(R0_out28),
.i0029(R0_in29),
.i0129(R0_out29),
.i0030(R0_in30),
.i0130(R0_out30),
.i0031(R0_in31),
.i0131(R0_out31),
.i0032(R0_in32),
.i0132(R0_out32),
.i0033(R0_in33),
.i0133(R0_out33),
.i0034(R0_in34),
.i0134(R0_out34),
.i0035(R0_in35),
.i0135(R0_out35),
.i0036(R0_in36),
.i0136(R0_out36),
.i0037(R0_in37),
.i0137(R0_out37),
.i0038(R0_in38),
.i0138(R0_out38),
.i0039(R0_in39),
.i0139(R0_out39),
.i0040(R0_in40),
.i0140(R0_out40),
.i0041(R0_in41),
.i0141(R0_out41),
.i0042(R0_in42),
.i0142(R0_out42),
.i0043(R0_in43),
.i0143(R0_out43),
.i0044(R0_in44),
.i0144(R0_out44),
.i0045(R0_in45),
.i0145(R0_out45),
.i0046(R0_in46),
.i0146(R0_out46),
.i0047(R0_in47),
.i0147(R0_out47),
.i0048(R0_in48),
.i0148(R0_out48),
.i0049(R0_in49),
.i0149(R0_out49),
.i0050(R0_in50),
.i0150(R0_out50),
.i0051(R0_in51),
.i0151(R0_out51),
.i0052(R0_in52),
.i0152(R0_out52),
.i0053(R0_in53),
.i0153(R0_out53),
.i0054(R0_in54),
.i0154(R0_out54),
.i0055(R0_in55),
.i0155(R0_out55),
.i0056(R0_in56),
.i0156(R0_out56),
.i0057(R0_in57),
.i0157(R0_out57),
.i0058(R0_in58),
.i0158(R0_out58),
.i0059(R0_in59),
.i0159(R0_out59),
.i0060(R0_in60),
.i0160(R0_out60),
.i0061(R0_in61),
.i0161(R0_out61),
.i0062(R0_in62),
.i0162(R0_out62)); //,
//.Write(Write),.Read(Read));
router r1
( .clk(clk), .rst(reset),
.i00(input_R0),
.i01(port1_inR0),
.o00(output_R0),
.o01(port1_outR0),.Write(Write),.Read(Read)
);
router r2
( .clk(clk), .rst(reset),
.i00(input_R1),
.i01(port1_inR1),
.o00(output_R1),
.o01(port1_outR1),.Write(Write),.Read(Read)
);
router r3
( .clk(clk), .rst(reset),
.i00(input_R2),
.i01(port1_inR2),
.o00(output_R2),
.o01(port1_outR2),.Write(Write),.Read(Read)
);
router r4
( .clk(clk), .rst(reset),
.i00(input_R3),
.i01(port1_inR3),
.o00(output_R3),
.o01(port1_outR3),.Write(Write),.Read(Read)
);
router r5
( .clk(clk), .rst(reset),
.i00(input_R4),
.i01(port1_inR4),
.o00(output_R4),
.o01(port1_outR4),.Write(Write),.Read(Read)
);
router r6
( .clk(clk), .rst(reset),
.i00(input_R5),
.i01(port1_inR5),
.o00(output_R5),
.o01(port1_outR5),.Write(Write),.Read(Read)
);
router r7
( .clk(clk), .rst(reset),
.i00(input_R6),
.i01(port1_inR6),
.o00(output_R6),
.o01(port1_outR6),.Write(Write),.Read(Read)
);
router r8
( .clk(clk), .rst(reset),
.i00(input_R7),
.i01(port1_inR7),
.o00(output_R7),
.o01(port1_outR7),.Write(Write),.Read(Read)
);
router r9
( .clk(clk), .rst(reset),
.i00(input_R8),
.i01(port1_inR8),
.o00(output_R8),
.o01(port1_outR8),.Write(Write),.Read(Read)
);
router r10
( .clk(clk), .rst(reset),
.i00(input_R9),
.i01(port1_inR9),
.o00(output_R9),
.o01(port1_outR9),.Write(Write),.Read(Read)
);
router r11
( .clk(clk), .rst(reset),
.i00(input_R10),
.i01(port1_inR10),
.o00(output_R10),
.o01(port1_outR10),.Write(Write),.Read(Read)
);
router r12
( .clk(clk), .rst(reset),
.i00(input_R11),
.i01(port1_inR11),
.o00(output_R11),
.o01(port1_outR11),.Write(Write),.Read(Read)
);
router r13
( .clk(clk), .rst(reset),
.i00(input_R12),
.i01(port1_inR12),
.o00(output_R12),
.o01(port1_outR12),.Write(Write),.Read(Read)
);
router r14
( .clk(clk), .rst(reset),
.i00(input_R13),
.i01(port1_inR13),
.o00(output_R13),
.o01(port1_outR13),.Write(Write),.Read(Read)
);
router r15
( .clk(clk), .rst(reset),
.i00(input_R14),
.i01(port1_inR14),
.o00(output_R14),
.o01(port1_outR14),.Write(Write),.Read(Read)
);
router r16
( .clk(clk), .rst(reset),
.i00(input_R15),
.i01(port1_inR15),
.o00(output_R15),
.o01(port1_outR15),.Write(Write),.Read(Read)
);
router r17
( .clk(clk), .rst(reset),
.i00(input_R16),
.i01(port1_inR16),
.o00(output_R16),
.o01(port1_outR16),.Write(Write),.Read(Read)
);
router r18
( .clk(clk), .rst(reset),
.i00(input_R17),
.i01(port1_inR17),
.o00(output_R17),
.o01(port1_outR17),.Write(Write),.Read(Read)
);
router r19
( .clk(clk), .rst(reset),
.i00(input_R18),
.i01(port1_inR18),
.o00(output_R18),
.o01(port1_outR18),.Write(Write),.Read(Read)
);
router r20
( .clk(clk), .rst(reset),
.i00(input_R19),
.i01(port1_inR19),
.o00(output_R19),
.o01(port1_outR19),.Write(Write),.Read(Read)
);
router r21
( .clk(clk), .rst(reset),
.i00(input_R20),
.i01(port1_inR20),
.o00(output_R20),
.o01(port1_outR20),.Write(Write),.Read(Read)
);
router r22
( .clk(clk), .rst(reset),
.i00(input_R21),
.i01(port1_inR21),
.o00(output_R21),
.o01(port1_outR21),.Write(Write),.Read(Read)
);
router r23
( .clk(clk), .rst(reset),
.i00(input_R22),
.i01(port1_inR22),
.o00(output_R22),
.o01(port1_outR22),.Write(Write),.Read(Read)
);
router r24
( .clk(clk), .rst(reset),
.i00(input_R23),
.i01(port1_inR23),
.o00(output_R23),
.o01(port1_outR23),.Write(Write),.Read(Read)
);
router r25
( .clk(clk), .rst(reset),
.i00(input_R24),
.i01(port1_inR24),
.o00(output_R24),
.o01(port1_outR24),.Write(Write),.Read(Read)
);
router r26
( .clk(clk), .rst(reset),
.i00(input_R25),
.i01(port1_inR25),
.o00(output_R25),
.o01(port1_outR25),.Write(Write),.Read(Read)
);
router r27
( .clk(clk), .rst(reset),
.i00(input_R26),
.i01(port1_inR26),
.o00(output_R26),
.o01(port1_outR26),.Write(Write),.Read(Read)
);
router r28
( .clk(clk), .rst(reset),
.i00(input_R27),
.i01(port1_inR27),
.o00(output_R27),
.o01(port1_outR27),.Write(Write),.Read(Read)
);
router r29
( .clk(clk), .rst(reset),
.i00(input_R28),
.i01(port1_inR28),
.o00(output_R28),
.o01(port1_outR28),.Write(Write),.Read(Read)
);
router r30
( .clk(clk), .rst(reset),
.i00(input_R29),
.i01(port1_inR29),
.o00(output_R29),
.o01(port1_outR29),.Write(Write),.Read(Read)
);
router r31
( .clk(clk), .rst(reset),
.i00(input_R30),
.i01(port1_inR30),
.o00(output_R30),
.o01(port1_outR30),.Write(Write),.Read(Read)
);
router r32
( .clk(clk), .rst(reset),
.i00(input_R31),
.i01(port1_inR31),
.o00(output_R31),
.o01(port1_outR31),.Write(Write),.Read(Read)
);
router r33
( .clk(clk), .rst(reset),
.i00(input_R32),
.i01(port1_inR32),
.o00(output_R32),
.o01(port1_outR32),.Write(Write),.Read(Read)
);
router r34
( .clk(clk), .rst(reset),
.i00(input_R33),
.i01(port1_inR33),
.o00(output_R33),
.o01(port1_outR33),.Write(Write),.Read(Read)
);
router r35
( .clk(clk), .rst(reset),
.i00(input_R34),
.i01(port1_inR34),
.o00(output_R34),
.o01(port1_outR34),.Write(Write),.Read(Read)
);
router r36
( .clk(clk), .rst(reset),
.i00(input_R35),
.i01(port1_inR35),
.o00(output_R35),
.o01(port1_outR35),.Write(Write),.Read(Read)
);
router r37
( .clk(clk), .rst(reset),
.i00(input_R36),
.i01(port1_inR36),
.o00(output_R36),
.o01(port1_outR36),.Write(Write),.Read(Read)
);
router r38
( .clk(clk), .rst(reset),
.i00(input_R37),
.i01(port1_inR37),
.o00(output_R37),
.o01(port1_outR37),.Write(Write),.Read(Read)
);
router r39
( .clk(clk), .rst(reset),
.i00(input_R38),
.i01(port1_inR38),
.o00(output_R38),
.o01(port1_outR38),.Write(Write),.Read(Read)
);
router r40
( .clk(clk), .rst(reset),
.i00(input_R39),
.i01(port1_inR39),
.o00(output_R39),
.o01(port1_outR39),.Write(Write),.Read(Read)
);
router r41
( .clk(clk), .rst(reset),
.i00(input_R40),
.i01(port1_inR40),
.o00(output_R40),
.o01(port1_outR40),.Write(Write),.Read(Read)
);
router r42
( .clk(clk), .rst(reset),
.i00(input_R41),
.i01(port1_inR41),
.o00(output_R41),
.o01(port1_outR41),.Write(Write),.Read(Read)
);
router r43
( .clk(clk), .rst(reset),
.i00(input_R42),
.i01(port1_inR42),
.o00(output_R42),
.o01(port1_outR42),.Write(Write),.Read(Read)
);
router r44
( .clk(clk), .rst(reset),
.i00(input_R43),
.i01(port1_inR43),
.o00(output_R43),
.o01(port1_outR43),.Write(Write),.Read(Read)
);
router r45
( .clk(clk), .rst(reset),
.i00(input_R44),
.i01(port1_inR44),
.o00(output_R44),
.o01(port1_outR44),.Write(Write),.Read(Read)
);
router r46
( .clk(clk), .rst(reset),
.i00(input_R45),
.i01(port1_inR45),
.o00(output_R45),
.o01(port1_outR45),.Write(Write),.Read(Read)
);
router r47
( .clk(clk), .rst(reset),
.i00(input_R46),
.i01(port1_inR46),
.o00(output_R46),
.o01(port1_outR46),.Write(Write),.Read(Read)
);
router r48
( .clk(clk), .rst(reset),
.i00(input_R47),
.i01(port1_inR47),
.o00(output_R47),
.o01(port1_outR47),.Write(Write),.Read(Read)
);
router r49
( .clk(clk), .rst(reset),
.i00(input_R48),
.i01(port1_inR48),
.o00(output_R48),
.o01(port1_outR48),.Write(Write),.Read(Read)
);
router r50
( .clk(clk), .rst(reset),
.i00(input_R49),
.i01(port1_inR49),
.o00(output_R49),
.o01(port1_outR49),.Write(Write),.Read(Read)
);
router r51
( .clk(clk), .rst(reset),
.i00(input_R50),
.i01(port1_inR50),
.o00(output_R50),
.o01(port1_outR50),.Write(Write),.Read(Read)
);
router r52
( .clk(clk), .rst(reset),
.i00(input_R51),
.i01(port1_inR51),
.o00(output_R51),
.o01(port1_outR51),.Write(Write),.Read(Read)
);
router r53
( .clk(clk), .rst(reset),
.i00(input_R52),
.i01(port1_inR52),
.o00(output_R52),
.o01(port1_outR52),.Write(Write),.Read(Read)
);
router r54
( .clk(clk), .rst(reset),
.i00(input_R53),
.i01(port1_inR53),
.o00(output_R53),
.o01(port1_outR53),.Write(Write),.Read(Read)
);
router r55
( .clk(clk), .rst(reset),
.i00(input_R54),
.i01(port1_inR54),
.o00(output_R54),
.o01(port1_outR54),.Write(Write),.Read(Read)
);
router r56
( .clk(clk), .rst(reset),
.i00(input_R55),
.i01(port1_inR55),
.o00(output_R55),
.o01(port1_outR55),.Write(Write),.Read(Read)
);
router r57
( .clk(clk), .rst(reset),
.i00(input_R56),
.i01(port1_inR56),
.o00(output_R56),
.o01(port1_outR56),.Write(Write),.Read(Read)
);
router r58
( .clk(clk), .rst(reset),
.i00(input_R57),
.i01(port1_inR57),
.o00(output_R57),
.o01(port1_outR57),.Write(Write),.Read(Read)
);
router r59
( .clk(clk), .rst(reset),
.i00(input_R58),
.i01(port1_inR58),
.o00(output_R58),
.o01(port1_outR58),.Write(Write),.Read(Read)
);
router r60
( .clk(clk), .rst(reset),
.i00(input_R59),
.i01(port1_inR59),
.o00(output_R59),
.o01(port1_outR59),.Write(Write),.Read(Read)
);
router r61
( .clk(clk), .rst(reset),
.i00(input_R60),
.i01(port1_inR60),
.o00(output_R60),
.o01(port1_outR60),.Write(Write),.Read(Read)
);
router r62
( .clk(clk), .rst(reset),
.i00(input_R61),
.i01(port1_inR61),
.o00(output_R61),
.o01(port1_outR61),.Write(Write),.Read(Read)
);
router r63
( .clk(clk), .rst(reset),
.i00(input_R62),
.i01(port1_inR62),
.o00(output_R62),
.o01(port1_outR62),.Write(Write),.Read(Read)
);
always @ ( posedge clk)
begin
port1_inR1<=R0_out0;
port1_inR2<=R0_out1;
port1_inR3<=R0_out2;
port1_inR4<=R0_out3;
port1_inR5<=R0_out4;
port1_inR6<=R0_out5;
port1_inR7<=R0_out6;
port1_inR8<=R0_out7;
port1_inR9<=R0_out8;
port1_inR10<=R0_out9;
port1_inR11<=R0_out10;
port1_inR12<=R0_out11;
port1_inR13<=R0_out12;
port1_inR14<=R0_out13;
port1_inR15<=R0_out14;
port1_inR16<=R0_out15;
port1_inR17<=R0_out16;
port1_inR18<=R0_out17;
port1_inR19<=R0_out18;
port1_inR20<=R0_out19;
port1_inR21<=R0_out20;
port1_inR22<=R0_out21;
port1_inR23<=R0_out22;
port1_inR24<=R0_out23;
port1_inR25<=R0_out24;
port1_inR26<=R0_out25;
port1_inR27<=R0_out26;
port1_inR28<=R0_out27;
port1_inR29<=R0_out28;
port1_inR30<=R0_out29;
port1_inR31<=R0_out30;
port1_inR32<=R0_out31;
port1_inR33<=R0_out32;
port1_inR34<=R0_out33;
port1_inR35<=R0_out34;
port1_inR36<=R0_out35;
port1_inR37<=R0_out36;
port1_inR38<=R0_out37;
port1_inR39<=R0_out38;
port1_inR40<=R0_out39;
port1_inR41<=R0_out40;
port1_inR42<=R0_out41;
port1_inR43<=R0_out42;
port1_inR44<=R0_out43;
port1_inR45<=R0_out44;
port1_inR46<=R0_out45;
port1_inR47<=R0_out46;
port1_inR48<=R0_out47;
port1_inR49<=R0_out48;
port1_inR50<=R0_out49;
port1_inR51<=R0_out50;
port1_inR52<=R0_out51;
port1_inR53<=R0_out52;
port1_inR54<=R0_out53;
port1_inR55<=R0_out54;
port1_inR56<=R0_out55;
port1_inR57<=R0_out56;
port1_inR58<=R0_out57;
port1_inR59<=R0_out58;
port1_inR60<=R0_out59;
port1_inR61<=R0_out60;
port1_inR62<=R0_out61;
port1_inR63<=R0_out62;
R0_in0<=port1_outR1;
R0_in1<=port1_outR2;
R0_in2<=port1_outR3;
R0_in3<=port1_outR4;
R0_in4<=port1_outR5;
R0_in5<=port1_outR6;
R0_in6<=port1_outR7;
R0_in7<=port1_outR8;
R0_in8<=port1_outR9;
R0_in9<=port1_outR10;
R0_in10<=port1_outR11;
R0_in11<=port1_outR12;
R0_in12<=port1_outR13;
R0_in13<=port1_outR14;
R0_in14<=port1_outR15;
R0_in15<=port1_outR16;
R0_in16<=port1_outR17;
R0_in17<=port1_outR18;
R0_in18<=port1_outR19;
R0_in19<=port1_outR20;
R0_in20<=port1_outR21;
R0_in21<=port1_outR22;
R0_in22<=port1_outR23;
R0_in23<=port1_outR24;
R0_in24<=port1_outR25;
R0_in25<=port1_outR26;
R0_in26<=port1_outR27;
R0_in27<=port1_outR28;
R0_in28<=port1_outR29;
R0_in29<=port1_outR30;
R0_in30<=port1_outR31;
R0_in31<=port1_outR32;
R0_in32<=port1_outR33;
R0_in33<=port1_outR34;
R0_in34<=port1_outR35;
R0_in35<=port1_outR36;
R0_in36<=port1_outR37;
R0_in37<=port1_outR38;
R0_in38<=port1_outR39;
R0_in39<=port1_outR40;
R0_in40<=port1_outR41;
R0_in41<=port1_outR42;
R0_in42<=port1_outR43;
R0_in43<=port1_outR44;
R0_in44<=port1_outR45;
R0_in45<=port1_outR46;
R0_in46<=port1_outR47;
R0_in47<=port1_outR48;
R0_in48<=port1_outR49;
R0_in49<=port1_outR50;
R0_in50<=port1_outR51;
R0_in51<=port1_outR52;
R0_in52<=port1_outR53;
R0_in53<=port1_outR54;
R0_in54<=port1_outR55;
R0_in55<=port1_outR56;
R0_in56<=port1_outR57;
R0_in57<=port1_outR58;
R0_in58<=port1_outR59;
R0_in59<=port1_outR60;
R0_in60<=port1_outR61;
R0_in61<=port1_outR62;
R0_in62<=port1_outR63;
end
endmodule
