module torus (
local0_in00,local0_out00,
local0_in01,local0_out01,
local0_in02,local0_out02,
local0_in03,local0_out03,
local0_in04,local0_out04,
local0_in05,local0_out05,
local0_in06,local0_out06,
local0_in07,local0_out07,
local0_in08,local0_out08,
local0_in09,local0_out09,
local0_in010,local0_out010,
local0_in011,local0_out011,
local0_in012,local0_out012,
local0_in013,local0_out013,
local0_in014,local0_out014,
local0_in015,local0_out015,
local1_in10,local1_out10,
local1_in11,local1_out11,
local1_in12,local1_out12,
local1_in13,local1_out13,
local1_in14,local1_out14,
local1_in15,local1_out15,
local1_in16,local1_out16,
local1_in17,local1_out17,
local1_in18,local1_out18,
local1_in19,local1_out19,
local1_in110,local1_out110,
local1_in111,local1_out111,
local1_in112,local1_out112,
local1_in113,local1_out113,
local1_in114,local1_out114,
local1_in115,local1_out115,
local2_in20,local2_out20,
local2_in21,local2_out21,
local2_in22,local2_out22,
local2_in23,local2_out23,
local2_in24,local2_out24,
local2_in25,local2_out25,
local2_in26,local2_out26,
local2_in27,local2_out27,
local2_in28,local2_out28,
local2_in29,local2_out29,
local2_in210,local2_out210,
local2_in211,local2_out211,
local2_in212,local2_out212,
local2_in213,local2_out213,
local2_in214,local2_out214,
local2_in215,local2_out215,
local3_in30,local3_out30,
local3_in31,local3_out31,
local3_in32,local3_out32,
local3_in33,local3_out33,
local3_in34,local3_out34,
local3_in35,local3_out35,
local3_in36,local3_out36,
local3_in37,local3_out37,
local3_in38,local3_out38,
local3_in39,local3_out39,
local3_in310,local3_out310,
local3_in311,local3_out311,
local3_in312,local3_out312,
local3_in313,local3_out313,
local3_in314,local3_out314,
local3_in315,local3_out315,
local4_in40,local4_out40,
local4_in41,local4_out41,
local4_in42,local4_out42,
local4_in43,local4_out43,
local4_in44,local4_out44,
local4_in45,local4_out45,
local4_in46,local4_out46,
local4_in47,local4_out47,
local4_in48,local4_out48,
local4_in49,local4_out49,
local4_in410,local4_out410,
local4_in411,local4_out411,
local4_in412,local4_out412,
local4_in413,local4_out413,
local4_in414,local4_out414,
local4_in415,local4_out415,
local5_in50,local5_out50,
local5_in51,local5_out51,
local5_in52,local5_out52,
local5_in53,local5_out53,
local5_in54,local5_out54,
local5_in55,local5_out55,
local5_in56,local5_out56,
local5_in57,local5_out57,
local5_in58,local5_out58,
local5_in59,local5_out59,
local5_in510,local5_out510,
local5_in511,local5_out511,
local5_in512,local5_out512,
local5_in513,local5_out513,
local5_in514,local5_out514,
local5_in515,local5_out515,
local6_in60,local6_out60,
local6_in61,local6_out61,
local6_in62,local6_out62,
local6_in63,local6_out63,
local6_in64,local6_out64,
local6_in65,local6_out65,
local6_in66,local6_out66,
local6_in67,local6_out67,
local6_in68,local6_out68,
local6_in69,local6_out69,
local6_in610,local6_out610,
local6_in611,local6_out611,
local6_in612,local6_out612,
local6_in613,local6_out613,
local6_in614,local6_out614,
local6_in615,local6_out615,
local7_in70,local7_out70,
local7_in71,local7_out71,
local7_in72,local7_out72,
local7_in73,local7_out73,
local7_in74,local7_out74,
local7_in75,local7_out75,
local7_in76,local7_out76,
local7_in77,local7_out77,
local7_in78,local7_out78,
local7_in79,local7_out79,
local7_in710,local7_out710,
local7_in711,local7_out711,
local7_in712,local7_out712,
local7_in713,local7_out713,
local7_in714,local7_out714,
local7_in715,local7_out715,
local8_in80,local8_out80,
local8_in81,local8_out81,
local8_in82,local8_out82,
local8_in83,local8_out83,
local8_in84,local8_out84,
local8_in85,local8_out85,
local8_in86,local8_out86,
local8_in87,local8_out87,
local8_in88,local8_out88,
local8_in89,local8_out89,
local8_in810,local8_out810,
local8_in811,local8_out811,
local8_in812,local8_out812,
local8_in813,local8_out813,
local8_in814,local8_out814,
local8_in815,local8_out815,
local9_in90,local9_out90,
local9_in91,local9_out91,
local9_in92,local9_out92,
local9_in93,local9_out93,
local9_in94,local9_out94,
local9_in95,local9_out95,
local9_in96,local9_out96,
local9_in97,local9_out97,
local9_in98,local9_out98,
local9_in99,local9_out99,
local9_in910,local9_out910,
local9_in911,local9_out911,
local9_in912,local9_out912,
local9_in913,local9_out913,
local9_in914,local9_out914,
local9_in915,local9_out915,
local10_in100,local10_out100,
local10_in101,local10_out101,
local10_in102,local10_out102,
local10_in103,local10_out103,
local10_in104,local10_out104,
local10_in105,local10_out105,
local10_in106,local10_out106,
local10_in107,local10_out107,
local10_in108,local10_out108,
local10_in109,local10_out109,
local10_in1010,local10_out1010,
local10_in1011,local10_out1011,
local10_in1012,local10_out1012,
local10_in1013,local10_out1013,
local10_in1014,local10_out1014,
local10_in1015,local10_out1015,
local11_in110,local11_out110,
local11_in111,local11_out111,
local11_in112,local11_out112,
local11_in113,local11_out113,
local11_in114,local11_out114,
local11_in115,local11_out115,
local11_in116,local11_out116,
local11_in117,local11_out117,
local11_in118,local11_out118,
local11_in119,local11_out119,
local11_in1110,local11_out1110,
local11_in1111,local11_out1111,
local11_in1112,local11_out1112,
local11_in1113,local11_out1113,
local11_in1114,local11_out1114,
local11_in1115,local11_out1115,
local12_in120,local12_out120,
local12_in121,local12_out121,
local12_in122,local12_out122,
local12_in123,local12_out123,
local12_in124,local12_out124,
local12_in125,local12_out125,
local12_in126,local12_out126,
local12_in127,local12_out127,
local12_in128,local12_out128,
local12_in129,local12_out129,
local12_in1210,local12_out1210,
local12_in1211,local12_out1211,
local12_in1212,local12_out1212,
local12_in1213,local12_out1213,
local12_in1214,local12_out1214,
local12_in1215,local12_out1215,
local13_in130,local13_out130,
local13_in131,local13_out131,
local13_in132,local13_out132,
local13_in133,local13_out133,
local13_in134,local13_out134,
local13_in135,local13_out135,
local13_in136,local13_out136,
local13_in137,local13_out137,
local13_in138,local13_out138,
local13_in139,local13_out139,
local13_in1310,local13_out1310,
local13_in1311,local13_out1311,
local13_in1312,local13_out1312,
local13_in1313,local13_out1313,
local13_in1314,local13_out1314,
local13_in1315,local13_out1315,
local14_in140,local14_out140,
local14_in141,local14_out141,
local14_in142,local14_out142,
local14_in143,local14_out143,
local14_in144,local14_out144,
local14_in145,local14_out145,
local14_in146,local14_out146,
local14_in147,local14_out147,
local14_in148,local14_out148,
local14_in149,local14_out149,
local14_in1410,local14_out1410,
local14_in1411,local14_out1411,
local14_in1412,local14_out1412,
local14_in1413,local14_out1413,
local14_in1414,local14_out1414,
local14_in1415,local14_out1415,
local15_in150,local15_out150,
local15_in151,local15_out151,
local15_in152,local15_out152,
local15_in153,local15_out153,
local15_in154,local15_out154,
local15_in155,local15_out155,
local15_in156,local15_out156,
local15_in157,local15_out157,
local15_in158,local15_out158,
local15_in159,local15_out159,
local15_in1510,local15_out1510,
local15_in1511,local15_out1511,
local15_in1512,local15_out1512,
local15_in1513,local15_out1513,
local15_in1514,local15_out1514,
local15_in1515,local15_out1515,
clk, reset,  Write, Read);
input clk, reset, Write, Read; 
parameter DATAWID = 32;
input [DATAWID-1:0] local0_in00;
output [DATAWID-1:0] local0_out00;
input [DATAWID-1:0] local0_in01;
output [DATAWID-1:0] local0_out01;
input [DATAWID-1:0] local0_in02;
output [DATAWID-1:0] local0_out02;
input [DATAWID-1:0] local0_in03;
output [DATAWID-1:0] local0_out03;
input [DATAWID-1:0] local0_in04;
output [DATAWID-1:0] local0_out04;
input [DATAWID-1:0] local0_in05;
output [DATAWID-1:0] local0_out05;
input [DATAWID-1:0] local0_in06;
output [DATAWID-1:0] local0_out06;
input [DATAWID-1:0] local0_in07;
output [DATAWID-1:0] local0_out07;
input [DATAWID-1:0] local0_in08;
output [DATAWID-1:0] local0_out08;
input [DATAWID-1:0] local0_in09;
output [DATAWID-1:0] local0_out09;
input [DATAWID-1:0] local0_in010;
output [DATAWID-1:0] local0_out010;
input [DATAWID-1:0] local0_in011;
output [DATAWID-1:0] local0_out011;
input [DATAWID-1:0] local0_in012;
output [DATAWID-1:0] local0_out012;
input [DATAWID-1:0] local0_in013;
output [DATAWID-1:0] local0_out013;
input [DATAWID-1:0] local0_in014;
output [DATAWID-1:0] local0_out014;
input [DATAWID-1:0] local0_in015;
output [DATAWID-1:0] local0_out015;
input [DATAWID-1:0] local1_in10;
output [DATAWID-1:0] local1_out10;
input [DATAWID-1:0] local1_in11;
output [DATAWID-1:0] local1_out11;
input [DATAWID-1:0] local1_in12;
output [DATAWID-1:0] local1_out12;
input [DATAWID-1:0] local1_in13;
output [DATAWID-1:0] local1_out13;
input [DATAWID-1:0] local1_in14;
output [DATAWID-1:0] local1_out14;
input [DATAWID-1:0] local1_in15;
output [DATAWID-1:0] local1_out15;
input [DATAWID-1:0] local1_in16;
output [DATAWID-1:0] local1_out16;
input [DATAWID-1:0] local1_in17;
output [DATAWID-1:0] local1_out17;
input [DATAWID-1:0] local1_in18;
output [DATAWID-1:0] local1_out18;
input [DATAWID-1:0] local1_in19;
output [DATAWID-1:0] local1_out19;
input [DATAWID-1:0] local1_in110;
output [DATAWID-1:0] local1_out110;
input [DATAWID-1:0] local1_in111;
output [DATAWID-1:0] local1_out111;
input [DATAWID-1:0] local1_in112;
output [DATAWID-1:0] local1_out112;
input [DATAWID-1:0] local1_in113;
output [DATAWID-1:0] local1_out113;
input [DATAWID-1:0] local1_in114;
output [DATAWID-1:0] local1_out114;
input [DATAWID-1:0] local1_in115;
output [DATAWID-1:0] local1_out115;
input [DATAWID-1:0] local2_in20;
output [DATAWID-1:0] local2_out20;
input [DATAWID-1:0] local2_in21;
output [DATAWID-1:0] local2_out21;
input [DATAWID-1:0] local2_in22;
output [DATAWID-1:0] local2_out22;
input [DATAWID-1:0] local2_in23;
output [DATAWID-1:0] local2_out23;
input [DATAWID-1:0] local2_in24;
output [DATAWID-1:0] local2_out24;
input [DATAWID-1:0] local2_in25;
output [DATAWID-1:0] local2_out25;
input [DATAWID-1:0] local2_in26;
output [DATAWID-1:0] local2_out26;
input [DATAWID-1:0] local2_in27;
output [DATAWID-1:0] local2_out27;
input [DATAWID-1:0] local2_in28;
output [DATAWID-1:0] local2_out28;
input [DATAWID-1:0] local2_in29;
output [DATAWID-1:0] local2_out29;
input [DATAWID-1:0] local2_in210;
output [DATAWID-1:0] local2_out210;
input [DATAWID-1:0] local2_in211;
output [DATAWID-1:0] local2_out211;
input [DATAWID-1:0] local2_in212;
output [DATAWID-1:0] local2_out212;
input [DATAWID-1:0] local2_in213;
output [DATAWID-1:0] local2_out213;
input [DATAWID-1:0] local2_in214;
output [DATAWID-1:0] local2_out214;
input [DATAWID-1:0] local2_in215;
output [DATAWID-1:0] local2_out215;
input [DATAWID-1:0] local3_in30;
output [DATAWID-1:0] local3_out30;
input [DATAWID-1:0] local3_in31;
output [DATAWID-1:0] local3_out31;
input [DATAWID-1:0] local3_in32;
output [DATAWID-1:0] local3_out32;
input [DATAWID-1:0] local3_in33;
output [DATAWID-1:0] local3_out33;
input [DATAWID-1:0] local3_in34;
output [DATAWID-1:0] local3_out34;
input [DATAWID-1:0] local3_in35;
output [DATAWID-1:0] local3_out35;
input [DATAWID-1:0] local3_in36;
output [DATAWID-1:0] local3_out36;
input [DATAWID-1:0] local3_in37;
output [DATAWID-1:0] local3_out37;
input [DATAWID-1:0] local3_in38;
output [DATAWID-1:0] local3_out38;
input [DATAWID-1:0] local3_in39;
output [DATAWID-1:0] local3_out39;
input [DATAWID-1:0] local3_in310;
output [DATAWID-1:0] local3_out310;
input [DATAWID-1:0] local3_in311;
output [DATAWID-1:0] local3_out311;
input [DATAWID-1:0] local3_in312;
output [DATAWID-1:0] local3_out312;
input [DATAWID-1:0] local3_in313;
output [DATAWID-1:0] local3_out313;
input [DATAWID-1:0] local3_in314;
output [DATAWID-1:0] local3_out314;
input [DATAWID-1:0] local3_in315;
output [DATAWID-1:0] local3_out315;
input [DATAWID-1:0] local4_in40;
output [DATAWID-1:0] local4_out40;
input [DATAWID-1:0] local4_in41;
output [DATAWID-1:0] local4_out41;
input [DATAWID-1:0] local4_in42;
output [DATAWID-1:0] local4_out42;
input [DATAWID-1:0] local4_in43;
output [DATAWID-1:0] local4_out43;
input [DATAWID-1:0] local4_in44;
output [DATAWID-1:0] local4_out44;
input [DATAWID-1:0] local4_in45;
output [DATAWID-1:0] local4_out45;
input [DATAWID-1:0] local4_in46;
output [DATAWID-1:0] local4_out46;
input [DATAWID-1:0] local4_in47;
output [DATAWID-1:0] local4_out47;
input [DATAWID-1:0] local4_in48;
output [DATAWID-1:0] local4_out48;
input [DATAWID-1:0] local4_in49;
output [DATAWID-1:0] local4_out49;
input [DATAWID-1:0] local4_in410;
output [DATAWID-1:0] local4_out410;
input [DATAWID-1:0] local4_in411;
output [DATAWID-1:0] local4_out411;
input [DATAWID-1:0] local4_in412;
output [DATAWID-1:0] local4_out412;
input [DATAWID-1:0] local4_in413;
output [DATAWID-1:0] local4_out413;
input [DATAWID-1:0] local4_in414;
output [DATAWID-1:0] local4_out414;
input [DATAWID-1:0] local4_in415;
output [DATAWID-1:0] local4_out415;
input [DATAWID-1:0] local5_in50;
output [DATAWID-1:0] local5_out50;
input [DATAWID-1:0] local5_in51;
output [DATAWID-1:0] local5_out51;
input [DATAWID-1:0] local5_in52;
output [DATAWID-1:0] local5_out52;
input [DATAWID-1:0] local5_in53;
output [DATAWID-1:0] local5_out53;
input [DATAWID-1:0] local5_in54;
output [DATAWID-1:0] local5_out54;
input [DATAWID-1:0] local5_in55;
output [DATAWID-1:0] local5_out55;
input [DATAWID-1:0] local5_in56;
output [DATAWID-1:0] local5_out56;
input [DATAWID-1:0] local5_in57;
output [DATAWID-1:0] local5_out57;
input [DATAWID-1:0] local5_in58;
output [DATAWID-1:0] local5_out58;
input [DATAWID-1:0] local5_in59;
output [DATAWID-1:0] local5_out59;
input [DATAWID-1:0] local5_in510;
output [DATAWID-1:0] local5_out510;
input [DATAWID-1:0] local5_in511;
output [DATAWID-1:0] local5_out511;
input [DATAWID-1:0] local5_in512;
output [DATAWID-1:0] local5_out512;
input [DATAWID-1:0] local5_in513;
output [DATAWID-1:0] local5_out513;
input [DATAWID-1:0] local5_in514;
output [DATAWID-1:0] local5_out514;
input [DATAWID-1:0] local5_in515;
output [DATAWID-1:0] local5_out515;
input [DATAWID-1:0] local6_in60;
output [DATAWID-1:0] local6_out60;
input [DATAWID-1:0] local6_in61;
output [DATAWID-1:0] local6_out61;
input [DATAWID-1:0] local6_in62;
output [DATAWID-1:0] local6_out62;
input [DATAWID-1:0] local6_in63;
output [DATAWID-1:0] local6_out63;
input [DATAWID-1:0] local6_in64;
output [DATAWID-1:0] local6_out64;
input [DATAWID-1:0] local6_in65;
output [DATAWID-1:0] local6_out65;
input [DATAWID-1:0] local6_in66;
output [DATAWID-1:0] local6_out66;
input [DATAWID-1:0] local6_in67;
output [DATAWID-1:0] local6_out67;
input [DATAWID-1:0] local6_in68;
output [DATAWID-1:0] local6_out68;
input [DATAWID-1:0] local6_in69;
output [DATAWID-1:0] local6_out69;
input [DATAWID-1:0] local6_in610;
output [DATAWID-1:0] local6_out610;
input [DATAWID-1:0] local6_in611;
output [DATAWID-1:0] local6_out611;
input [DATAWID-1:0] local6_in612;
output [DATAWID-1:0] local6_out612;
input [DATAWID-1:0] local6_in613;
output [DATAWID-1:0] local6_out613;
input [DATAWID-1:0] local6_in614;
output [DATAWID-1:0] local6_out614;
input [DATAWID-1:0] local6_in615;
output [DATAWID-1:0] local6_out615;
input [DATAWID-1:0] local7_in70;
output [DATAWID-1:0] local7_out70;
input [DATAWID-1:0] local7_in71;
output [DATAWID-1:0] local7_out71;
input [DATAWID-1:0] local7_in72;
output [DATAWID-1:0] local7_out72;
input [DATAWID-1:0] local7_in73;
output [DATAWID-1:0] local7_out73;
input [DATAWID-1:0] local7_in74;
output [DATAWID-1:0] local7_out74;
input [DATAWID-1:0] local7_in75;
output [DATAWID-1:0] local7_out75;
input [DATAWID-1:0] local7_in76;
output [DATAWID-1:0] local7_out76;
input [DATAWID-1:0] local7_in77;
output [DATAWID-1:0] local7_out77;
input [DATAWID-1:0] local7_in78;
output [DATAWID-1:0] local7_out78;
input [DATAWID-1:0] local7_in79;
output [DATAWID-1:0] local7_out79;
input [DATAWID-1:0] local7_in710;
output [DATAWID-1:0] local7_out710;
input [DATAWID-1:0] local7_in711;
output [DATAWID-1:0] local7_out711;
input [DATAWID-1:0] local7_in712;
output [DATAWID-1:0] local7_out712;
input [DATAWID-1:0] local7_in713;
output [DATAWID-1:0] local7_out713;
input [DATAWID-1:0] local7_in714;
output [DATAWID-1:0] local7_out714;
input [DATAWID-1:0] local7_in715;
output [DATAWID-1:0] local7_out715;
input [DATAWID-1:0] local8_in80;
output [DATAWID-1:0] local8_out80;
input [DATAWID-1:0] local8_in81;
output [DATAWID-1:0] local8_out81;
input [DATAWID-1:0] local8_in82;
output [DATAWID-1:0] local8_out82;
input [DATAWID-1:0] local8_in83;
output [DATAWID-1:0] local8_out83;
input [DATAWID-1:0] local8_in84;
output [DATAWID-1:0] local8_out84;
input [DATAWID-1:0] local8_in85;
output [DATAWID-1:0] local8_out85;
input [DATAWID-1:0] local8_in86;
output [DATAWID-1:0] local8_out86;
input [DATAWID-1:0] local8_in87;
output [DATAWID-1:0] local8_out87;
input [DATAWID-1:0] local8_in88;
output [DATAWID-1:0] local8_out88;
input [DATAWID-1:0] local8_in89;
output [DATAWID-1:0] local8_out89;
input [DATAWID-1:0] local8_in810;
output [DATAWID-1:0] local8_out810;
input [DATAWID-1:0] local8_in811;
output [DATAWID-1:0] local8_out811;
input [DATAWID-1:0] local8_in812;
output [DATAWID-1:0] local8_out812;
input [DATAWID-1:0] local8_in813;
output [DATAWID-1:0] local8_out813;
input [DATAWID-1:0] local8_in814;
output [DATAWID-1:0] local8_out814;
input [DATAWID-1:0] local8_in815;
output [DATAWID-1:0] local8_out815;
input [DATAWID-1:0] local9_in90;
output [DATAWID-1:0] local9_out90;
input [DATAWID-1:0] local9_in91;
output [DATAWID-1:0] local9_out91;
input [DATAWID-1:0] local9_in92;
output [DATAWID-1:0] local9_out92;
input [DATAWID-1:0] local9_in93;
output [DATAWID-1:0] local9_out93;
input [DATAWID-1:0] local9_in94;
output [DATAWID-1:0] local9_out94;
input [DATAWID-1:0] local9_in95;
output [DATAWID-1:0] local9_out95;
input [DATAWID-1:0] local9_in96;
output [DATAWID-1:0] local9_out96;
input [DATAWID-1:0] local9_in97;
output [DATAWID-1:0] local9_out97;
input [DATAWID-1:0] local9_in98;
output [DATAWID-1:0] local9_out98;
input [DATAWID-1:0] local9_in99;
output [DATAWID-1:0] local9_out99;
input [DATAWID-1:0] local9_in910;
output [DATAWID-1:0] local9_out910;
input [DATAWID-1:0] local9_in911;
output [DATAWID-1:0] local9_out911;
input [DATAWID-1:0] local9_in912;
output [DATAWID-1:0] local9_out912;
input [DATAWID-1:0] local9_in913;
output [DATAWID-1:0] local9_out913;
input [DATAWID-1:0] local9_in914;
output [DATAWID-1:0] local9_out914;
input [DATAWID-1:0] local9_in915;
output [DATAWID-1:0] local9_out915;
input [DATAWID-1:0] local10_in100;
output [DATAWID-1:0] local10_out100;
input [DATAWID-1:0] local10_in101;
output [DATAWID-1:0] local10_out101;
input [DATAWID-1:0] local10_in102;
output [DATAWID-1:0] local10_out102;
input [DATAWID-1:0] local10_in103;
output [DATAWID-1:0] local10_out103;
input [DATAWID-1:0] local10_in104;
output [DATAWID-1:0] local10_out104;
input [DATAWID-1:0] local10_in105;
output [DATAWID-1:0] local10_out105;
input [DATAWID-1:0] local10_in106;
output [DATAWID-1:0] local10_out106;
input [DATAWID-1:0] local10_in107;
output [DATAWID-1:0] local10_out107;
input [DATAWID-1:0] local10_in108;
output [DATAWID-1:0] local10_out108;
input [DATAWID-1:0] local10_in109;
output [DATAWID-1:0] local10_out109;
input [DATAWID-1:0] local10_in1010;
output [DATAWID-1:0] local10_out1010;
input [DATAWID-1:0] local10_in1011;
output [DATAWID-1:0] local10_out1011;
input [DATAWID-1:0] local10_in1012;
output [DATAWID-1:0] local10_out1012;
input [DATAWID-1:0] local10_in1013;
output [DATAWID-1:0] local10_out1013;
input [DATAWID-1:0] local10_in1014;
output [DATAWID-1:0] local10_out1014;
input [DATAWID-1:0] local10_in1015;
output [DATAWID-1:0] local10_out1015;
input [DATAWID-1:0] local11_in110;
output [DATAWID-1:0] local11_out110;
input [DATAWID-1:0] local11_in111;
output [DATAWID-1:0] local11_out111;
input [DATAWID-1:0] local11_in112;
output [DATAWID-1:0] local11_out112;
input [DATAWID-1:0] local11_in113;
output [DATAWID-1:0] local11_out113;
input [DATAWID-1:0] local11_in114;
output [DATAWID-1:0] local11_out114;
input [DATAWID-1:0] local11_in115;
output [DATAWID-1:0] local11_out115;
input [DATAWID-1:0] local11_in116;
output [DATAWID-1:0] local11_out116;
input [DATAWID-1:0] local11_in117;
output [DATAWID-1:0] local11_out117;
input [DATAWID-1:0] local11_in118;
output [DATAWID-1:0] local11_out118;
input [DATAWID-1:0] local11_in119;
output [DATAWID-1:0] local11_out119;
input [DATAWID-1:0] local11_in1110;
output [DATAWID-1:0] local11_out1110;
input [DATAWID-1:0] local11_in1111;
output [DATAWID-1:0] local11_out1111;
input [DATAWID-1:0] local11_in1112;
output [DATAWID-1:0] local11_out1112;
input [DATAWID-1:0] local11_in1113;
output [DATAWID-1:0] local11_out1113;
input [DATAWID-1:0] local11_in1114;
output [DATAWID-1:0] local11_out1114;
input [DATAWID-1:0] local11_in1115;
output [DATAWID-1:0] local11_out1115;
input [DATAWID-1:0] local12_in120;
output [DATAWID-1:0] local12_out120;
input [DATAWID-1:0] local12_in121;
output [DATAWID-1:0] local12_out121;
input [DATAWID-1:0] local12_in122;
output [DATAWID-1:0] local12_out122;
input [DATAWID-1:0] local12_in123;
output [DATAWID-1:0] local12_out123;
input [DATAWID-1:0] local12_in124;
output [DATAWID-1:0] local12_out124;
input [DATAWID-1:0] local12_in125;
output [DATAWID-1:0] local12_out125;
input [DATAWID-1:0] local12_in126;
output [DATAWID-1:0] local12_out126;
input [DATAWID-1:0] local12_in127;
output [DATAWID-1:0] local12_out127;
input [DATAWID-1:0] local12_in128;
output [DATAWID-1:0] local12_out128;
input [DATAWID-1:0] local12_in129;
output [DATAWID-1:0] local12_out129;
input [DATAWID-1:0] local12_in1210;
output [DATAWID-1:0] local12_out1210;
input [DATAWID-1:0] local12_in1211;
output [DATAWID-1:0] local12_out1211;
input [DATAWID-1:0] local12_in1212;
output [DATAWID-1:0] local12_out1212;
input [DATAWID-1:0] local12_in1213;
output [DATAWID-1:0] local12_out1213;
input [DATAWID-1:0] local12_in1214;
output [DATAWID-1:0] local12_out1214;
input [DATAWID-1:0] local12_in1215;
output [DATAWID-1:0] local12_out1215;
input [DATAWID-1:0] local13_in130;
output [DATAWID-1:0] local13_out130;
input [DATAWID-1:0] local13_in131;
output [DATAWID-1:0] local13_out131;
input [DATAWID-1:0] local13_in132;
output [DATAWID-1:0] local13_out132;
input [DATAWID-1:0] local13_in133;
output [DATAWID-1:0] local13_out133;
input [DATAWID-1:0] local13_in134;
output [DATAWID-1:0] local13_out134;
input [DATAWID-1:0] local13_in135;
output [DATAWID-1:0] local13_out135;
input [DATAWID-1:0] local13_in136;
output [DATAWID-1:0] local13_out136;
input [DATAWID-1:0] local13_in137;
output [DATAWID-1:0] local13_out137;
input [DATAWID-1:0] local13_in138;
output [DATAWID-1:0] local13_out138;
input [DATAWID-1:0] local13_in139;
output [DATAWID-1:0] local13_out139;
input [DATAWID-1:0] local13_in1310;
output [DATAWID-1:0] local13_out1310;
input [DATAWID-1:0] local13_in1311;
output [DATAWID-1:0] local13_out1311;
input [DATAWID-1:0] local13_in1312;
output [DATAWID-1:0] local13_out1312;
input [DATAWID-1:0] local13_in1313;
output [DATAWID-1:0] local13_out1313;
input [DATAWID-1:0] local13_in1314;
output [DATAWID-1:0] local13_out1314;
input [DATAWID-1:0] local13_in1315;
output [DATAWID-1:0] local13_out1315;
input [DATAWID-1:0] local14_in140;
output [DATAWID-1:0] local14_out140;
input [DATAWID-1:0] local14_in141;
output [DATAWID-1:0] local14_out141;
input [DATAWID-1:0] local14_in142;
output [DATAWID-1:0] local14_out142;
input [DATAWID-1:0] local14_in143;
output [DATAWID-1:0] local14_out143;
input [DATAWID-1:0] local14_in144;
output [DATAWID-1:0] local14_out144;
input [DATAWID-1:0] local14_in145;
output [DATAWID-1:0] local14_out145;
input [DATAWID-1:0] local14_in146;
output [DATAWID-1:0] local14_out146;
input [DATAWID-1:0] local14_in147;
output [DATAWID-1:0] local14_out147;
input [DATAWID-1:0] local14_in148;
output [DATAWID-1:0] local14_out148;
input [DATAWID-1:0] local14_in149;
output [DATAWID-1:0] local14_out149;
input [DATAWID-1:0] local14_in1410;
output [DATAWID-1:0] local14_out1410;
input [DATAWID-1:0] local14_in1411;
output [DATAWID-1:0] local14_out1411;
input [DATAWID-1:0] local14_in1412;
output [DATAWID-1:0] local14_out1412;
input [DATAWID-1:0] local14_in1413;
output [DATAWID-1:0] local14_out1413;
input [DATAWID-1:0] local14_in1414;
output [DATAWID-1:0] local14_out1414;
input [DATAWID-1:0] local14_in1415;
output [DATAWID-1:0] local14_out1415;
input [DATAWID-1:0] local15_in150;
output [DATAWID-1:0] local15_out150;
input [DATAWID-1:0] local15_in151;
output [DATAWID-1:0] local15_out151;
input [DATAWID-1:0] local15_in152;
output [DATAWID-1:0] local15_out152;
input [DATAWID-1:0] local15_in153;
output [DATAWID-1:0] local15_out153;
input [DATAWID-1:0] local15_in154;
output [DATAWID-1:0] local15_out154;
input [DATAWID-1:0] local15_in155;
output [DATAWID-1:0] local15_out155;
input [DATAWID-1:0] local15_in156;
output [DATAWID-1:0] local15_out156;
input [DATAWID-1:0] local15_in157;
output [DATAWID-1:0] local15_out157;
input [DATAWID-1:0] local15_in158;
output [DATAWID-1:0] local15_out158;
input [DATAWID-1:0] local15_in159;
output [DATAWID-1:0] local15_out159;
input [DATAWID-1:0] local15_in1510;
output [DATAWID-1:0] local15_out1510;
input [DATAWID-1:0] local15_in1511;
output [DATAWID-1:0] local15_out1511;
input [DATAWID-1:0] local15_in1512;
output [DATAWID-1:0] local15_out1512;
input [DATAWID-1:0] local15_in1513;
output [DATAWID-1:0] local15_out1513;
input [DATAWID-1:0] local15_in1514;
output [DATAWID-1:0] local15_out1514;
input [DATAWID-1:0] local15_in1515;
output [DATAWID-1:0] local15_out1515;
reg [DATAWID-1:0] east0_in00;
reg [DATAWID-1:0] west0_in00;
reg [DATAWID-1:0] north0_in00;
reg [DATAWID-1:0] south0_in00;
reg [DATAWID-1:0] east0_in01;
reg [DATAWID-1:0] west0_in01;
reg [DATAWID-1:0] north0_in01;
reg [DATAWID-1:0] south0_in01;
reg [DATAWID-1:0] east0_in02;
reg [DATAWID-1:0] west0_in02;
reg [DATAWID-1:0] north0_in02;
reg [DATAWID-1:0] south0_in02;
reg [DATAWID-1:0] east0_in03;
reg [DATAWID-1:0] west0_in03;
reg [DATAWID-1:0] north0_in03;
reg [DATAWID-1:0] south0_in03;
reg [DATAWID-1:0] east0_in04;
reg [DATAWID-1:0] west0_in04;
reg [DATAWID-1:0] north0_in04;
reg [DATAWID-1:0] south0_in04;
reg [DATAWID-1:0] east0_in05;
reg [DATAWID-1:0] west0_in05;
reg [DATAWID-1:0] north0_in05;
reg [DATAWID-1:0] south0_in05;
reg [DATAWID-1:0] east0_in06;
reg [DATAWID-1:0] west0_in06;
reg [DATAWID-1:0] north0_in06;
reg [DATAWID-1:0] south0_in06;
reg [DATAWID-1:0] east0_in07;
reg [DATAWID-1:0] west0_in07;
reg [DATAWID-1:0] north0_in07;
reg [DATAWID-1:0] south0_in07;
reg [DATAWID-1:0] east0_in08;
reg [DATAWID-1:0] west0_in08;
reg [DATAWID-1:0] north0_in08;
reg [DATAWID-1:0] south0_in08;
reg [DATAWID-1:0] east0_in09;
reg [DATAWID-1:0] west0_in09;
reg [DATAWID-1:0] north0_in09;
reg [DATAWID-1:0] south0_in09;
reg [DATAWID-1:0] east0_in010;
reg [DATAWID-1:0] west0_in010;
reg [DATAWID-1:0] north0_in010;
reg [DATAWID-1:0] south0_in010;
reg [DATAWID-1:0] east0_in011;
reg [DATAWID-1:0] west0_in011;
reg [DATAWID-1:0] north0_in011;
reg [DATAWID-1:0] south0_in011;
reg [DATAWID-1:0] east0_in012;
reg [DATAWID-1:0] west0_in012;
reg [DATAWID-1:0] north0_in012;
reg [DATAWID-1:0] south0_in012;
reg [DATAWID-1:0] east0_in013;
reg [DATAWID-1:0] west0_in013;
reg [DATAWID-1:0] north0_in013;
reg [DATAWID-1:0] south0_in013;
reg [DATAWID-1:0] east0_in014;
reg [DATAWID-1:0] west0_in014;
reg [DATAWID-1:0] north0_in014;
reg [DATAWID-1:0] south0_in014;
reg [DATAWID-1:0] east0_in015;
reg [DATAWID-1:0] west0_in015;
reg [DATAWID-1:0] north0_in015;
reg [DATAWID-1:0] south0_in015;
reg [DATAWID-1:0] east1_in10;
reg [DATAWID-1:0] west1_in10;
reg [DATAWID-1:0] north1_in10;
reg [DATAWID-1:0] south1_in10;
reg [DATAWID-1:0] east1_in11;
reg [DATAWID-1:0] west1_in11;
reg [DATAWID-1:0] north1_in11;
reg [DATAWID-1:0] south1_in11;
reg [DATAWID-1:0] east1_in12;
reg [DATAWID-1:0] west1_in12;
reg [DATAWID-1:0] north1_in12;
reg [DATAWID-1:0] south1_in12;
reg [DATAWID-1:0] east1_in13;
reg [DATAWID-1:0] west1_in13;
reg [DATAWID-1:0] north1_in13;
reg [DATAWID-1:0] south1_in13;
reg [DATAWID-1:0] east1_in14;
reg [DATAWID-1:0] west1_in14;
reg [DATAWID-1:0] north1_in14;
reg [DATAWID-1:0] south1_in14;
reg [DATAWID-1:0] east1_in15;
reg [DATAWID-1:0] west1_in15;
reg [DATAWID-1:0] north1_in15;
reg [DATAWID-1:0] south1_in15;
reg [DATAWID-1:0] east1_in16;
reg [DATAWID-1:0] west1_in16;
reg [DATAWID-1:0] north1_in16;
reg [DATAWID-1:0] south1_in16;
reg [DATAWID-1:0] east1_in17;
reg [DATAWID-1:0] west1_in17;
reg [DATAWID-1:0] north1_in17;
reg [DATAWID-1:0] south1_in17;
reg [DATAWID-1:0] east1_in18;
reg [DATAWID-1:0] west1_in18;
reg [DATAWID-1:0] north1_in18;
reg [DATAWID-1:0] south1_in18;
reg [DATAWID-1:0] east1_in19;
reg [DATAWID-1:0] west1_in19;
reg [DATAWID-1:0] north1_in19;
reg [DATAWID-1:0] south1_in19;
reg [DATAWID-1:0] east1_in110;
reg [DATAWID-1:0] west1_in110;
reg [DATAWID-1:0] north1_in110;
reg [DATAWID-1:0] south1_in110;
reg [DATAWID-1:0] east1_in111;
reg [DATAWID-1:0] west1_in111;
reg [DATAWID-1:0] north1_in111;
reg [DATAWID-1:0] south1_in111;
reg [DATAWID-1:0] east1_in112;
reg [DATAWID-1:0] west1_in112;
reg [DATAWID-1:0] north1_in112;
reg [DATAWID-1:0] south1_in112;
reg [DATAWID-1:0] east1_in113;
reg [DATAWID-1:0] west1_in113;
reg [DATAWID-1:0] north1_in113;
reg [DATAWID-1:0] south1_in113;
reg [DATAWID-1:0] east1_in114;
reg [DATAWID-1:0] west1_in114;
reg [DATAWID-1:0] north1_in114;
reg [DATAWID-1:0] south1_in114;
reg [DATAWID-1:0] east1_in115;
reg [DATAWID-1:0] west1_in115;
reg [DATAWID-1:0] north1_in115;
reg [DATAWID-1:0] south1_in115;
reg [DATAWID-1:0] east2_in20;
reg [DATAWID-1:0] west2_in20;
reg [DATAWID-1:0] north2_in20;
reg [DATAWID-1:0] south2_in20;
reg [DATAWID-1:0] east2_in21;
reg [DATAWID-1:0] west2_in21;
reg [DATAWID-1:0] north2_in21;
reg [DATAWID-1:0] south2_in21;
reg [DATAWID-1:0] east2_in22;
reg [DATAWID-1:0] west2_in22;
reg [DATAWID-1:0] north2_in22;
reg [DATAWID-1:0] south2_in22;
reg [DATAWID-1:0] east2_in23;
reg [DATAWID-1:0] west2_in23;
reg [DATAWID-1:0] north2_in23;
reg [DATAWID-1:0] south2_in23;
reg [DATAWID-1:0] east2_in24;
reg [DATAWID-1:0] west2_in24;
reg [DATAWID-1:0] north2_in24;
reg [DATAWID-1:0] south2_in24;
reg [DATAWID-1:0] east2_in25;
reg [DATAWID-1:0] west2_in25;
reg [DATAWID-1:0] north2_in25;
reg [DATAWID-1:0] south2_in25;
reg [DATAWID-1:0] east2_in26;
reg [DATAWID-1:0] west2_in26;
reg [DATAWID-1:0] north2_in26;
reg [DATAWID-1:0] south2_in26;
reg [DATAWID-1:0] east2_in27;
reg [DATAWID-1:0] west2_in27;
reg [DATAWID-1:0] north2_in27;
reg [DATAWID-1:0] south2_in27;
reg [DATAWID-1:0] east2_in28;
reg [DATAWID-1:0] west2_in28;
reg [DATAWID-1:0] north2_in28;
reg [DATAWID-1:0] south2_in28;
reg [DATAWID-1:0] east2_in29;
reg [DATAWID-1:0] west2_in29;
reg [DATAWID-1:0] north2_in29;
reg [DATAWID-1:0] south2_in29;
reg [DATAWID-1:0] east2_in210;
reg [DATAWID-1:0] west2_in210;
reg [DATAWID-1:0] north2_in210;
reg [DATAWID-1:0] south2_in210;
reg [DATAWID-1:0] east2_in211;
reg [DATAWID-1:0] west2_in211;
reg [DATAWID-1:0] north2_in211;
reg [DATAWID-1:0] south2_in211;
reg [DATAWID-1:0] east2_in212;
reg [DATAWID-1:0] west2_in212;
reg [DATAWID-1:0] north2_in212;
reg [DATAWID-1:0] south2_in212;
reg [DATAWID-1:0] east2_in213;
reg [DATAWID-1:0] west2_in213;
reg [DATAWID-1:0] north2_in213;
reg [DATAWID-1:0] south2_in213;
reg [DATAWID-1:0] east2_in214;
reg [DATAWID-1:0] west2_in214;
reg [DATAWID-1:0] north2_in214;
reg [DATAWID-1:0] south2_in214;
reg [DATAWID-1:0] east2_in215;
reg [DATAWID-1:0] west2_in215;
reg [DATAWID-1:0] north2_in215;
reg [DATAWID-1:0] south2_in215;
reg [DATAWID-1:0] east3_in30;
reg [DATAWID-1:0] west3_in30;
reg [DATAWID-1:0] north3_in30;
reg [DATAWID-1:0] south3_in30;
reg [DATAWID-1:0] east3_in31;
reg [DATAWID-1:0] west3_in31;
reg [DATAWID-1:0] north3_in31;
reg [DATAWID-1:0] south3_in31;
reg [DATAWID-1:0] east3_in32;
reg [DATAWID-1:0] west3_in32;
reg [DATAWID-1:0] north3_in32;
reg [DATAWID-1:0] south3_in32;
reg [DATAWID-1:0] east3_in33;
reg [DATAWID-1:0] west3_in33;
reg [DATAWID-1:0] north3_in33;
reg [DATAWID-1:0] south3_in33;
reg [DATAWID-1:0] east3_in34;
reg [DATAWID-1:0] west3_in34;
reg [DATAWID-1:0] north3_in34;
reg [DATAWID-1:0] south3_in34;
reg [DATAWID-1:0] east3_in35;
reg [DATAWID-1:0] west3_in35;
reg [DATAWID-1:0] north3_in35;
reg [DATAWID-1:0] south3_in35;
reg [DATAWID-1:0] east3_in36;
reg [DATAWID-1:0] west3_in36;
reg [DATAWID-1:0] north3_in36;
reg [DATAWID-1:0] south3_in36;
reg [DATAWID-1:0] east3_in37;
reg [DATAWID-1:0] west3_in37;
reg [DATAWID-1:0] north3_in37;
reg [DATAWID-1:0] south3_in37;
reg [DATAWID-1:0] east3_in38;
reg [DATAWID-1:0] west3_in38;
reg [DATAWID-1:0] north3_in38;
reg [DATAWID-1:0] south3_in38;
reg [DATAWID-1:0] east3_in39;
reg [DATAWID-1:0] west3_in39;
reg [DATAWID-1:0] north3_in39;
reg [DATAWID-1:0] south3_in39;
reg [DATAWID-1:0] east3_in310;
reg [DATAWID-1:0] west3_in310;
reg [DATAWID-1:0] north3_in310;
reg [DATAWID-1:0] south3_in310;
reg [DATAWID-1:0] east3_in311;
reg [DATAWID-1:0] west3_in311;
reg [DATAWID-1:0] north3_in311;
reg [DATAWID-1:0] south3_in311;
reg [DATAWID-1:0] east3_in312;
reg [DATAWID-1:0] west3_in312;
reg [DATAWID-1:0] north3_in312;
reg [DATAWID-1:0] south3_in312;
reg [DATAWID-1:0] east3_in313;
reg [DATAWID-1:0] west3_in313;
reg [DATAWID-1:0] north3_in313;
reg [DATAWID-1:0] south3_in313;
reg [DATAWID-1:0] east3_in314;
reg [DATAWID-1:0] west3_in314;
reg [DATAWID-1:0] north3_in314;
reg [DATAWID-1:0] south3_in314;
reg [DATAWID-1:0] east3_in315;
reg [DATAWID-1:0] west3_in315;
reg [DATAWID-1:0] north3_in315;
reg [DATAWID-1:0] south3_in315;
reg [DATAWID-1:0] east4_in40;
reg [DATAWID-1:0] west4_in40;
reg [DATAWID-1:0] north4_in40;
reg [DATAWID-1:0] south4_in40;
reg [DATAWID-1:0] east4_in41;
reg [DATAWID-1:0] west4_in41;
reg [DATAWID-1:0] north4_in41;
reg [DATAWID-1:0] south4_in41;
reg [DATAWID-1:0] east4_in42;
reg [DATAWID-1:0] west4_in42;
reg [DATAWID-1:0] north4_in42;
reg [DATAWID-1:0] south4_in42;
reg [DATAWID-1:0] east4_in43;
reg [DATAWID-1:0] west4_in43;
reg [DATAWID-1:0] north4_in43;
reg [DATAWID-1:0] south4_in43;
reg [DATAWID-1:0] east4_in44;
reg [DATAWID-1:0] west4_in44;
reg [DATAWID-1:0] north4_in44;
reg [DATAWID-1:0] south4_in44;
reg [DATAWID-1:0] east4_in45;
reg [DATAWID-1:0] west4_in45;
reg [DATAWID-1:0] north4_in45;
reg [DATAWID-1:0] south4_in45;
reg [DATAWID-1:0] east4_in46;
reg [DATAWID-1:0] west4_in46;
reg [DATAWID-1:0] north4_in46;
reg [DATAWID-1:0] south4_in46;
reg [DATAWID-1:0] east4_in47;
reg [DATAWID-1:0] west4_in47;
reg [DATAWID-1:0] north4_in47;
reg [DATAWID-1:0] south4_in47;
reg [DATAWID-1:0] east4_in48;
reg [DATAWID-1:0] west4_in48;
reg [DATAWID-1:0] north4_in48;
reg [DATAWID-1:0] south4_in48;
reg [DATAWID-1:0] east4_in49;
reg [DATAWID-1:0] west4_in49;
reg [DATAWID-1:0] north4_in49;
reg [DATAWID-1:0] south4_in49;
reg [DATAWID-1:0] east4_in410;
reg [DATAWID-1:0] west4_in410;
reg [DATAWID-1:0] north4_in410;
reg [DATAWID-1:0] south4_in410;
reg [DATAWID-1:0] east4_in411;
reg [DATAWID-1:0] west4_in411;
reg [DATAWID-1:0] north4_in411;
reg [DATAWID-1:0] south4_in411;
reg [DATAWID-1:0] east4_in412;
reg [DATAWID-1:0] west4_in412;
reg [DATAWID-1:0] north4_in412;
reg [DATAWID-1:0] south4_in412;
reg [DATAWID-1:0] east4_in413;
reg [DATAWID-1:0] west4_in413;
reg [DATAWID-1:0] north4_in413;
reg [DATAWID-1:0] south4_in413;
reg [DATAWID-1:0] east4_in414;
reg [DATAWID-1:0] west4_in414;
reg [DATAWID-1:0] north4_in414;
reg [DATAWID-1:0] south4_in414;
reg [DATAWID-1:0] east4_in415;
reg [DATAWID-1:0] west4_in415;
reg [DATAWID-1:0] north4_in415;
reg [DATAWID-1:0] south4_in415;
reg [DATAWID-1:0] east5_in50;
reg [DATAWID-1:0] west5_in50;
reg [DATAWID-1:0] north5_in50;
reg [DATAWID-1:0] south5_in50;
reg [DATAWID-1:0] east5_in51;
reg [DATAWID-1:0] west5_in51;
reg [DATAWID-1:0] north5_in51;
reg [DATAWID-1:0] south5_in51;
reg [DATAWID-1:0] east5_in52;
reg [DATAWID-1:0] west5_in52;
reg [DATAWID-1:0] north5_in52;
reg [DATAWID-1:0] south5_in52;
reg [DATAWID-1:0] east5_in53;
reg [DATAWID-1:0] west5_in53;
reg [DATAWID-1:0] north5_in53;
reg [DATAWID-1:0] south5_in53;
reg [DATAWID-1:0] east5_in54;
reg [DATAWID-1:0] west5_in54;
reg [DATAWID-1:0] north5_in54;
reg [DATAWID-1:0] south5_in54;
reg [DATAWID-1:0] east5_in55;
reg [DATAWID-1:0] west5_in55;
reg [DATAWID-1:0] north5_in55;
reg [DATAWID-1:0] south5_in55;
reg [DATAWID-1:0] east5_in56;
reg [DATAWID-1:0] west5_in56;
reg [DATAWID-1:0] north5_in56;
reg [DATAWID-1:0] south5_in56;
reg [DATAWID-1:0] east5_in57;
reg [DATAWID-1:0] west5_in57;
reg [DATAWID-1:0] north5_in57;
reg [DATAWID-1:0] south5_in57;
reg [DATAWID-1:0] east5_in58;
reg [DATAWID-1:0] west5_in58;
reg [DATAWID-1:0] north5_in58;
reg [DATAWID-1:0] south5_in58;
reg [DATAWID-1:0] east5_in59;
reg [DATAWID-1:0] west5_in59;
reg [DATAWID-1:0] north5_in59;
reg [DATAWID-1:0] south5_in59;
reg [DATAWID-1:0] east5_in510;
reg [DATAWID-1:0] west5_in510;
reg [DATAWID-1:0] north5_in510;
reg [DATAWID-1:0] south5_in510;
reg [DATAWID-1:0] east5_in511;
reg [DATAWID-1:0] west5_in511;
reg [DATAWID-1:0] north5_in511;
reg [DATAWID-1:0] south5_in511;
reg [DATAWID-1:0] east5_in512;
reg [DATAWID-1:0] west5_in512;
reg [DATAWID-1:0] north5_in512;
reg [DATAWID-1:0] south5_in512;
reg [DATAWID-1:0] east5_in513;
reg [DATAWID-1:0] west5_in513;
reg [DATAWID-1:0] north5_in513;
reg [DATAWID-1:0] south5_in513;
reg [DATAWID-1:0] east5_in514;
reg [DATAWID-1:0] west5_in514;
reg [DATAWID-1:0] north5_in514;
reg [DATAWID-1:0] south5_in514;
reg [DATAWID-1:0] east5_in515;
reg [DATAWID-1:0] west5_in515;
reg [DATAWID-1:0] north5_in515;
reg [DATAWID-1:0] south5_in515;
reg [DATAWID-1:0] east6_in60;
reg [DATAWID-1:0] west6_in60;
reg [DATAWID-1:0] north6_in60;
reg [DATAWID-1:0] south6_in60;
reg [DATAWID-1:0] east6_in61;
reg [DATAWID-1:0] west6_in61;
reg [DATAWID-1:0] north6_in61;
reg [DATAWID-1:0] south6_in61;
reg [DATAWID-1:0] east6_in62;
reg [DATAWID-1:0] west6_in62;
reg [DATAWID-1:0] north6_in62;
reg [DATAWID-1:0] south6_in62;
reg [DATAWID-1:0] east6_in63;
reg [DATAWID-1:0] west6_in63;
reg [DATAWID-1:0] north6_in63;
reg [DATAWID-1:0] south6_in63;
reg [DATAWID-1:0] east6_in64;
reg [DATAWID-1:0] west6_in64;
reg [DATAWID-1:0] north6_in64;
reg [DATAWID-1:0] south6_in64;
reg [DATAWID-1:0] east6_in65;
reg [DATAWID-1:0] west6_in65;
reg [DATAWID-1:0] north6_in65;
reg [DATAWID-1:0] south6_in65;
reg [DATAWID-1:0] east6_in66;
reg [DATAWID-1:0] west6_in66;
reg [DATAWID-1:0] north6_in66;
reg [DATAWID-1:0] south6_in66;
reg [DATAWID-1:0] east6_in67;
reg [DATAWID-1:0] west6_in67;
reg [DATAWID-1:0] north6_in67;
reg [DATAWID-1:0] south6_in67;
reg [DATAWID-1:0] east6_in68;
reg [DATAWID-1:0] west6_in68;
reg [DATAWID-1:0] north6_in68;
reg [DATAWID-1:0] south6_in68;
reg [DATAWID-1:0] east6_in69;
reg [DATAWID-1:0] west6_in69;
reg [DATAWID-1:0] north6_in69;
reg [DATAWID-1:0] south6_in69;
reg [DATAWID-1:0] east6_in610;
reg [DATAWID-1:0] west6_in610;
reg [DATAWID-1:0] north6_in610;
reg [DATAWID-1:0] south6_in610;
reg [DATAWID-1:0] east6_in611;
reg [DATAWID-1:0] west6_in611;
reg [DATAWID-1:0] north6_in611;
reg [DATAWID-1:0] south6_in611;
reg [DATAWID-1:0] east6_in612;
reg [DATAWID-1:0] west6_in612;
reg [DATAWID-1:0] north6_in612;
reg [DATAWID-1:0] south6_in612;
reg [DATAWID-1:0] east6_in613;
reg [DATAWID-1:0] west6_in613;
reg [DATAWID-1:0] north6_in613;
reg [DATAWID-1:0] south6_in613;
reg [DATAWID-1:0] east6_in614;
reg [DATAWID-1:0] west6_in614;
reg [DATAWID-1:0] north6_in614;
reg [DATAWID-1:0] south6_in614;
reg [DATAWID-1:0] east6_in615;
reg [DATAWID-1:0] west6_in615;
reg [DATAWID-1:0] north6_in615;
reg [DATAWID-1:0] south6_in615;
reg [DATAWID-1:0] east7_in70;
reg [DATAWID-1:0] west7_in70;
reg [DATAWID-1:0] north7_in70;
reg [DATAWID-1:0] south7_in70;
reg [DATAWID-1:0] east7_in71;
reg [DATAWID-1:0] west7_in71;
reg [DATAWID-1:0] north7_in71;
reg [DATAWID-1:0] south7_in71;
reg [DATAWID-1:0] east7_in72;
reg [DATAWID-1:0] west7_in72;
reg [DATAWID-1:0] north7_in72;
reg [DATAWID-1:0] south7_in72;
reg [DATAWID-1:0] east7_in73;
reg [DATAWID-1:0] west7_in73;
reg [DATAWID-1:0] north7_in73;
reg [DATAWID-1:0] south7_in73;
reg [DATAWID-1:0] east7_in74;
reg [DATAWID-1:0] west7_in74;
reg [DATAWID-1:0] north7_in74;
reg [DATAWID-1:0] south7_in74;
reg [DATAWID-1:0] east7_in75;
reg [DATAWID-1:0] west7_in75;
reg [DATAWID-1:0] north7_in75;
reg [DATAWID-1:0] south7_in75;
reg [DATAWID-1:0] east7_in76;
reg [DATAWID-1:0] west7_in76;
reg [DATAWID-1:0] north7_in76;
reg [DATAWID-1:0] south7_in76;
reg [DATAWID-1:0] east7_in77;
reg [DATAWID-1:0] west7_in77;
reg [DATAWID-1:0] north7_in77;
reg [DATAWID-1:0] south7_in77;
reg [DATAWID-1:0] east7_in78;
reg [DATAWID-1:0] west7_in78;
reg [DATAWID-1:0] north7_in78;
reg [DATAWID-1:0] south7_in78;
reg [DATAWID-1:0] east7_in79;
reg [DATAWID-1:0] west7_in79;
reg [DATAWID-1:0] north7_in79;
reg [DATAWID-1:0] south7_in79;
reg [DATAWID-1:0] east7_in710;
reg [DATAWID-1:0] west7_in710;
reg [DATAWID-1:0] north7_in710;
reg [DATAWID-1:0] south7_in710;
reg [DATAWID-1:0] east7_in711;
reg [DATAWID-1:0] west7_in711;
reg [DATAWID-1:0] north7_in711;
reg [DATAWID-1:0] south7_in711;
reg [DATAWID-1:0] east7_in712;
reg [DATAWID-1:0] west7_in712;
reg [DATAWID-1:0] north7_in712;
reg [DATAWID-1:0] south7_in712;
reg [DATAWID-1:0] east7_in713;
reg [DATAWID-1:0] west7_in713;
reg [DATAWID-1:0] north7_in713;
reg [DATAWID-1:0] south7_in713;
reg [DATAWID-1:0] east7_in714;
reg [DATAWID-1:0] west7_in714;
reg [DATAWID-1:0] north7_in714;
reg [DATAWID-1:0] south7_in714;
reg [DATAWID-1:0] east7_in715;
reg [DATAWID-1:0] west7_in715;
reg [DATAWID-1:0] north7_in715;
reg [DATAWID-1:0] south7_in715;
reg [DATAWID-1:0] east8_in80;
reg [DATAWID-1:0] west8_in80;
reg [DATAWID-1:0] north8_in80;
reg [DATAWID-1:0] south8_in80;
reg [DATAWID-1:0] east8_in81;
reg [DATAWID-1:0] west8_in81;
reg [DATAWID-1:0] north8_in81;
reg [DATAWID-1:0] south8_in81;
reg [DATAWID-1:0] east8_in82;
reg [DATAWID-1:0] west8_in82;
reg [DATAWID-1:0] north8_in82;
reg [DATAWID-1:0] south8_in82;
reg [DATAWID-1:0] east8_in83;
reg [DATAWID-1:0] west8_in83;
reg [DATAWID-1:0] north8_in83;
reg [DATAWID-1:0] south8_in83;
reg [DATAWID-1:0] east8_in84;
reg [DATAWID-1:0] west8_in84;
reg [DATAWID-1:0] north8_in84;
reg [DATAWID-1:0] south8_in84;
reg [DATAWID-1:0] east8_in85;
reg [DATAWID-1:0] west8_in85;
reg [DATAWID-1:0] north8_in85;
reg [DATAWID-1:0] south8_in85;
reg [DATAWID-1:0] east8_in86;
reg [DATAWID-1:0] west8_in86;
reg [DATAWID-1:0] north8_in86;
reg [DATAWID-1:0] south8_in86;
reg [DATAWID-1:0] east8_in87;
reg [DATAWID-1:0] west8_in87;
reg [DATAWID-1:0] north8_in87;
reg [DATAWID-1:0] south8_in87;
reg [DATAWID-1:0] east8_in88;
reg [DATAWID-1:0] west8_in88;
reg [DATAWID-1:0] north8_in88;
reg [DATAWID-1:0] south8_in88;
reg [DATAWID-1:0] east8_in89;
reg [DATAWID-1:0] west8_in89;
reg [DATAWID-1:0] north8_in89;
reg [DATAWID-1:0] south8_in89;
reg [DATAWID-1:0] east8_in810;
reg [DATAWID-1:0] west8_in810;
reg [DATAWID-1:0] north8_in810;
reg [DATAWID-1:0] south8_in810;
reg [DATAWID-1:0] east8_in811;
reg [DATAWID-1:0] west8_in811;
reg [DATAWID-1:0] north8_in811;
reg [DATAWID-1:0] south8_in811;
reg [DATAWID-1:0] east8_in812;
reg [DATAWID-1:0] west8_in812;
reg [DATAWID-1:0] north8_in812;
reg [DATAWID-1:0] south8_in812;
reg [DATAWID-1:0] east8_in813;
reg [DATAWID-1:0] west8_in813;
reg [DATAWID-1:0] north8_in813;
reg [DATAWID-1:0] south8_in813;
reg [DATAWID-1:0] east8_in814;
reg [DATAWID-1:0] west8_in814;
reg [DATAWID-1:0] north8_in814;
reg [DATAWID-1:0] south8_in814;
reg [DATAWID-1:0] east8_in815;
reg [DATAWID-1:0] west8_in815;
reg [DATAWID-1:0] north8_in815;
reg [DATAWID-1:0] south8_in815;
reg [DATAWID-1:0] east9_in90;
reg [DATAWID-1:0] west9_in90;
reg [DATAWID-1:0] north9_in90;
reg [DATAWID-1:0] south9_in90;
reg [DATAWID-1:0] east9_in91;
reg [DATAWID-1:0] west9_in91;
reg [DATAWID-1:0] north9_in91;
reg [DATAWID-1:0] south9_in91;
reg [DATAWID-1:0] east9_in92;
reg [DATAWID-1:0] west9_in92;
reg [DATAWID-1:0] north9_in92;
reg [DATAWID-1:0] south9_in92;
reg [DATAWID-1:0] east9_in93;
reg [DATAWID-1:0] west9_in93;
reg [DATAWID-1:0] north9_in93;
reg [DATAWID-1:0] south9_in93;
reg [DATAWID-1:0] east9_in94;
reg [DATAWID-1:0] west9_in94;
reg [DATAWID-1:0] north9_in94;
reg [DATAWID-1:0] south9_in94;
reg [DATAWID-1:0] east9_in95;
reg [DATAWID-1:0] west9_in95;
reg [DATAWID-1:0] north9_in95;
reg [DATAWID-1:0] south9_in95;
reg [DATAWID-1:0] east9_in96;
reg [DATAWID-1:0] west9_in96;
reg [DATAWID-1:0] north9_in96;
reg [DATAWID-1:0] south9_in96;
reg [DATAWID-1:0] east9_in97;
reg [DATAWID-1:0] west9_in97;
reg [DATAWID-1:0] north9_in97;
reg [DATAWID-1:0] south9_in97;
reg [DATAWID-1:0] east9_in98;
reg [DATAWID-1:0] west9_in98;
reg [DATAWID-1:0] north9_in98;
reg [DATAWID-1:0] south9_in98;
reg [DATAWID-1:0] east9_in99;
reg [DATAWID-1:0] west9_in99;
reg [DATAWID-1:0] north9_in99;
reg [DATAWID-1:0] south9_in99;
reg [DATAWID-1:0] east9_in910;
reg [DATAWID-1:0] west9_in910;
reg [DATAWID-1:0] north9_in910;
reg [DATAWID-1:0] south9_in910;
reg [DATAWID-1:0] east9_in911;
reg [DATAWID-1:0] west9_in911;
reg [DATAWID-1:0] north9_in911;
reg [DATAWID-1:0] south9_in911;
reg [DATAWID-1:0] east9_in912;
reg [DATAWID-1:0] west9_in912;
reg [DATAWID-1:0] north9_in912;
reg [DATAWID-1:0] south9_in912;
reg [DATAWID-1:0] east9_in913;
reg [DATAWID-1:0] west9_in913;
reg [DATAWID-1:0] north9_in913;
reg [DATAWID-1:0] south9_in913;
reg [DATAWID-1:0] east9_in914;
reg [DATAWID-1:0] west9_in914;
reg [DATAWID-1:0] north9_in914;
reg [DATAWID-1:0] south9_in914;
reg [DATAWID-1:0] east9_in915;
reg [DATAWID-1:0] west9_in915;
reg [DATAWID-1:0] north9_in915;
reg [DATAWID-1:0] south9_in915;
reg [DATAWID-1:0] east10_in100;
reg [DATAWID-1:0] west10_in100;
reg [DATAWID-1:0] north10_in100;
reg [DATAWID-1:0] south10_in100;
reg [DATAWID-1:0] east10_in101;
reg [DATAWID-1:0] west10_in101;
reg [DATAWID-1:0] north10_in101;
reg [DATAWID-1:0] south10_in101;
reg [DATAWID-1:0] east10_in102;
reg [DATAWID-1:0] west10_in102;
reg [DATAWID-1:0] north10_in102;
reg [DATAWID-1:0] south10_in102;
reg [DATAWID-1:0] east10_in103;
reg [DATAWID-1:0] west10_in103;
reg [DATAWID-1:0] north10_in103;
reg [DATAWID-1:0] south10_in103;
reg [DATAWID-1:0] east10_in104;
reg [DATAWID-1:0] west10_in104;
reg [DATAWID-1:0] north10_in104;
reg [DATAWID-1:0] south10_in104;
reg [DATAWID-1:0] east10_in105;
reg [DATAWID-1:0] west10_in105;
reg [DATAWID-1:0] north10_in105;
reg [DATAWID-1:0] south10_in105;
reg [DATAWID-1:0] east10_in106;
reg [DATAWID-1:0] west10_in106;
reg [DATAWID-1:0] north10_in106;
reg [DATAWID-1:0] south10_in106;
reg [DATAWID-1:0] east10_in107;
reg [DATAWID-1:0] west10_in107;
reg [DATAWID-1:0] north10_in107;
reg [DATAWID-1:0] south10_in107;
reg [DATAWID-1:0] east10_in108;
reg [DATAWID-1:0] west10_in108;
reg [DATAWID-1:0] north10_in108;
reg [DATAWID-1:0] south10_in108;
reg [DATAWID-1:0] east10_in109;
reg [DATAWID-1:0] west10_in109;
reg [DATAWID-1:0] north10_in109;
reg [DATAWID-1:0] south10_in109;
reg [DATAWID-1:0] east10_in1010;
reg [DATAWID-1:0] west10_in1010;
reg [DATAWID-1:0] north10_in1010;
reg [DATAWID-1:0] south10_in1010;
reg [DATAWID-1:0] east10_in1011;
reg [DATAWID-1:0] west10_in1011;
reg [DATAWID-1:0] north10_in1011;
reg [DATAWID-1:0] south10_in1011;
reg [DATAWID-1:0] east10_in1012;
reg [DATAWID-1:0] west10_in1012;
reg [DATAWID-1:0] north10_in1012;
reg [DATAWID-1:0] south10_in1012;
reg [DATAWID-1:0] east10_in1013;
reg [DATAWID-1:0] west10_in1013;
reg [DATAWID-1:0] north10_in1013;
reg [DATAWID-1:0] south10_in1013;
reg [DATAWID-1:0] east10_in1014;
reg [DATAWID-1:0] west10_in1014;
reg [DATAWID-1:0] north10_in1014;
reg [DATAWID-1:0] south10_in1014;
reg [DATAWID-1:0] east10_in1015;
reg [DATAWID-1:0] west10_in1015;
reg [DATAWID-1:0] north10_in1015;
reg [DATAWID-1:0] south10_in1015;
reg [DATAWID-1:0] east11_in110;
reg [DATAWID-1:0] west11_in110;
reg [DATAWID-1:0] north11_in110;
reg [DATAWID-1:0] south11_in110;
reg [DATAWID-1:0] east11_in111;
reg [DATAWID-1:0] west11_in111;
reg [DATAWID-1:0] north11_in111;
reg [DATAWID-1:0] south11_in111;
reg [DATAWID-1:0] east11_in112;
reg [DATAWID-1:0] west11_in112;
reg [DATAWID-1:0] north11_in112;
reg [DATAWID-1:0] south11_in112;
reg [DATAWID-1:0] east11_in113;
reg [DATAWID-1:0] west11_in113;
reg [DATAWID-1:0] north11_in113;
reg [DATAWID-1:0] south11_in113;
reg [DATAWID-1:0] east11_in114;
reg [DATAWID-1:0] west11_in114;
reg [DATAWID-1:0] north11_in114;
reg [DATAWID-1:0] south11_in114;
reg [DATAWID-1:0] east11_in115;
reg [DATAWID-1:0] west11_in115;
reg [DATAWID-1:0] north11_in115;
reg [DATAWID-1:0] south11_in115;
reg [DATAWID-1:0] east11_in116;
reg [DATAWID-1:0] west11_in116;
reg [DATAWID-1:0] north11_in116;
reg [DATAWID-1:0] south11_in116;
reg [DATAWID-1:0] east11_in117;
reg [DATAWID-1:0] west11_in117;
reg [DATAWID-1:0] north11_in117;
reg [DATAWID-1:0] south11_in117;
reg [DATAWID-1:0] east11_in118;
reg [DATAWID-1:0] west11_in118;
reg [DATAWID-1:0] north11_in118;
reg [DATAWID-1:0] south11_in118;
reg [DATAWID-1:0] east11_in119;
reg [DATAWID-1:0] west11_in119;
reg [DATAWID-1:0] north11_in119;
reg [DATAWID-1:0] south11_in119;
reg [DATAWID-1:0] east11_in1110;
reg [DATAWID-1:0] west11_in1110;
reg [DATAWID-1:0] north11_in1110;
reg [DATAWID-1:0] south11_in1110;
reg [DATAWID-1:0] east11_in1111;
reg [DATAWID-1:0] west11_in1111;
reg [DATAWID-1:0] north11_in1111;
reg [DATAWID-1:0] south11_in1111;
reg [DATAWID-1:0] east11_in1112;
reg [DATAWID-1:0] west11_in1112;
reg [DATAWID-1:0] north11_in1112;
reg [DATAWID-1:0] south11_in1112;
reg [DATAWID-1:0] east11_in1113;
reg [DATAWID-1:0] west11_in1113;
reg [DATAWID-1:0] north11_in1113;
reg [DATAWID-1:0] south11_in1113;
reg [DATAWID-1:0] east11_in1114;
reg [DATAWID-1:0] west11_in1114;
reg [DATAWID-1:0] north11_in1114;
reg [DATAWID-1:0] south11_in1114;
reg [DATAWID-1:0] east11_in1115;
reg [DATAWID-1:0] west11_in1115;
reg [DATAWID-1:0] north11_in1115;
reg [DATAWID-1:0] south11_in1115;
reg [DATAWID-1:0] east12_in120;
reg [DATAWID-1:0] west12_in120;
reg [DATAWID-1:0] north12_in120;
reg [DATAWID-1:0] south12_in120;
reg [DATAWID-1:0] east12_in121;
reg [DATAWID-1:0] west12_in121;
reg [DATAWID-1:0] north12_in121;
reg [DATAWID-1:0] south12_in121;
reg [DATAWID-1:0] east12_in122;
reg [DATAWID-1:0] west12_in122;
reg [DATAWID-1:0] north12_in122;
reg [DATAWID-1:0] south12_in122;
reg [DATAWID-1:0] east12_in123;
reg [DATAWID-1:0] west12_in123;
reg [DATAWID-1:0] north12_in123;
reg [DATAWID-1:0] south12_in123;
reg [DATAWID-1:0] east12_in124;
reg [DATAWID-1:0] west12_in124;
reg [DATAWID-1:0] north12_in124;
reg [DATAWID-1:0] south12_in124;
reg [DATAWID-1:0] east12_in125;
reg [DATAWID-1:0] west12_in125;
reg [DATAWID-1:0] north12_in125;
reg [DATAWID-1:0] south12_in125;
reg [DATAWID-1:0] east12_in126;
reg [DATAWID-1:0] west12_in126;
reg [DATAWID-1:0] north12_in126;
reg [DATAWID-1:0] south12_in126;
reg [DATAWID-1:0] east12_in127;
reg [DATAWID-1:0] west12_in127;
reg [DATAWID-1:0] north12_in127;
reg [DATAWID-1:0] south12_in127;
reg [DATAWID-1:0] east12_in128;
reg [DATAWID-1:0] west12_in128;
reg [DATAWID-1:0] north12_in128;
reg [DATAWID-1:0] south12_in128;
reg [DATAWID-1:0] east12_in129;
reg [DATAWID-1:0] west12_in129;
reg [DATAWID-1:0] north12_in129;
reg [DATAWID-1:0] south12_in129;
reg [DATAWID-1:0] east12_in1210;
reg [DATAWID-1:0] west12_in1210;
reg [DATAWID-1:0] north12_in1210;
reg [DATAWID-1:0] south12_in1210;
reg [DATAWID-1:0] east12_in1211;
reg [DATAWID-1:0] west12_in1211;
reg [DATAWID-1:0] north12_in1211;
reg [DATAWID-1:0] south12_in1211;
reg [DATAWID-1:0] east12_in1212;
reg [DATAWID-1:0] west12_in1212;
reg [DATAWID-1:0] north12_in1212;
reg [DATAWID-1:0] south12_in1212;
reg [DATAWID-1:0] east12_in1213;
reg [DATAWID-1:0] west12_in1213;
reg [DATAWID-1:0] north12_in1213;
reg [DATAWID-1:0] south12_in1213;
reg [DATAWID-1:0] east12_in1214;
reg [DATAWID-1:0] west12_in1214;
reg [DATAWID-1:0] north12_in1214;
reg [DATAWID-1:0] south12_in1214;
reg [DATAWID-1:0] east12_in1215;
reg [DATAWID-1:0] west12_in1215;
reg [DATAWID-1:0] north12_in1215;
reg [DATAWID-1:0] south12_in1215;
reg [DATAWID-1:0] east13_in130;
reg [DATAWID-1:0] west13_in130;
reg [DATAWID-1:0] north13_in130;
reg [DATAWID-1:0] south13_in130;
reg [DATAWID-1:0] east13_in131;
reg [DATAWID-1:0] west13_in131;
reg [DATAWID-1:0] north13_in131;
reg [DATAWID-1:0] south13_in131;
reg [DATAWID-1:0] east13_in132;
reg [DATAWID-1:0] west13_in132;
reg [DATAWID-1:0] north13_in132;
reg [DATAWID-1:0] south13_in132;
reg [DATAWID-1:0] east13_in133;
reg [DATAWID-1:0] west13_in133;
reg [DATAWID-1:0] north13_in133;
reg [DATAWID-1:0] south13_in133;
reg [DATAWID-1:0] east13_in134;
reg [DATAWID-1:0] west13_in134;
reg [DATAWID-1:0] north13_in134;
reg [DATAWID-1:0] south13_in134;
reg [DATAWID-1:0] east13_in135;
reg [DATAWID-1:0] west13_in135;
reg [DATAWID-1:0] north13_in135;
reg [DATAWID-1:0] south13_in135;
reg [DATAWID-1:0] east13_in136;
reg [DATAWID-1:0] west13_in136;
reg [DATAWID-1:0] north13_in136;
reg [DATAWID-1:0] south13_in136;
reg [DATAWID-1:0] east13_in137;
reg [DATAWID-1:0] west13_in137;
reg [DATAWID-1:0] north13_in137;
reg [DATAWID-1:0] south13_in137;
reg [DATAWID-1:0] east13_in138;
reg [DATAWID-1:0] west13_in138;
reg [DATAWID-1:0] north13_in138;
reg [DATAWID-1:0] south13_in138;
reg [DATAWID-1:0] east13_in139;
reg [DATAWID-1:0] west13_in139;
reg [DATAWID-1:0] north13_in139;
reg [DATAWID-1:0] south13_in139;
reg [DATAWID-1:0] east13_in1310;
reg [DATAWID-1:0] west13_in1310;
reg [DATAWID-1:0] north13_in1310;
reg [DATAWID-1:0] south13_in1310;
reg [DATAWID-1:0] east13_in1311;
reg [DATAWID-1:0] west13_in1311;
reg [DATAWID-1:0] north13_in1311;
reg [DATAWID-1:0] south13_in1311;
reg [DATAWID-1:0] east13_in1312;
reg [DATAWID-1:0] west13_in1312;
reg [DATAWID-1:0] north13_in1312;
reg [DATAWID-1:0] south13_in1312;
reg [DATAWID-1:0] east13_in1313;
reg [DATAWID-1:0] west13_in1313;
reg [DATAWID-1:0] north13_in1313;
reg [DATAWID-1:0] south13_in1313;
reg [DATAWID-1:0] east13_in1314;
reg [DATAWID-1:0] west13_in1314;
reg [DATAWID-1:0] north13_in1314;
reg [DATAWID-1:0] south13_in1314;
reg [DATAWID-1:0] east13_in1315;
reg [DATAWID-1:0] west13_in1315;
reg [DATAWID-1:0] north13_in1315;
reg [DATAWID-1:0] south13_in1315;
reg [DATAWID-1:0] east14_in140;
reg [DATAWID-1:0] west14_in140;
reg [DATAWID-1:0] north14_in140;
reg [DATAWID-1:0] south14_in140;
reg [DATAWID-1:0] east14_in141;
reg [DATAWID-1:0] west14_in141;
reg [DATAWID-1:0] north14_in141;
reg [DATAWID-1:0] south14_in141;
reg [DATAWID-1:0] east14_in142;
reg [DATAWID-1:0] west14_in142;
reg [DATAWID-1:0] north14_in142;
reg [DATAWID-1:0] south14_in142;
reg [DATAWID-1:0] east14_in143;
reg [DATAWID-1:0] west14_in143;
reg [DATAWID-1:0] north14_in143;
reg [DATAWID-1:0] south14_in143;
reg [DATAWID-1:0] east14_in144;
reg [DATAWID-1:0] west14_in144;
reg [DATAWID-1:0] north14_in144;
reg [DATAWID-1:0] south14_in144;
reg [DATAWID-1:0] east14_in145;
reg [DATAWID-1:0] west14_in145;
reg [DATAWID-1:0] north14_in145;
reg [DATAWID-1:0] south14_in145;
reg [DATAWID-1:0] east14_in146;
reg [DATAWID-1:0] west14_in146;
reg [DATAWID-1:0] north14_in146;
reg [DATAWID-1:0] south14_in146;
reg [DATAWID-1:0] east14_in147;
reg [DATAWID-1:0] west14_in147;
reg [DATAWID-1:0] north14_in147;
reg [DATAWID-1:0] south14_in147;
reg [DATAWID-1:0] east14_in148;
reg [DATAWID-1:0] west14_in148;
reg [DATAWID-1:0] north14_in148;
reg [DATAWID-1:0] south14_in148;
reg [DATAWID-1:0] east14_in149;
reg [DATAWID-1:0] west14_in149;
reg [DATAWID-1:0] north14_in149;
reg [DATAWID-1:0] south14_in149;
reg [DATAWID-1:0] east14_in1410;
reg [DATAWID-1:0] west14_in1410;
reg [DATAWID-1:0] north14_in1410;
reg [DATAWID-1:0] south14_in1410;
reg [DATAWID-1:0] east14_in1411;
reg [DATAWID-1:0] west14_in1411;
reg [DATAWID-1:0] north14_in1411;
reg [DATAWID-1:0] south14_in1411;
reg [DATAWID-1:0] east14_in1412;
reg [DATAWID-1:0] west14_in1412;
reg [DATAWID-1:0] north14_in1412;
reg [DATAWID-1:0] south14_in1412;
reg [DATAWID-1:0] east14_in1413;
reg [DATAWID-1:0] west14_in1413;
reg [DATAWID-1:0] north14_in1413;
reg [DATAWID-1:0] south14_in1413;
reg [DATAWID-1:0] east14_in1414;
reg [DATAWID-1:0] west14_in1414;
reg [DATAWID-1:0] north14_in1414;
reg [DATAWID-1:0] south14_in1414;
reg [DATAWID-1:0] east14_in1415;
reg [DATAWID-1:0] west14_in1415;
reg [DATAWID-1:0] north14_in1415;
reg [DATAWID-1:0] south14_in1415;
reg [DATAWID-1:0] east15_in150;
reg [DATAWID-1:0] west15_in150;
reg [DATAWID-1:0] north15_in150;
reg [DATAWID-1:0] south15_in150;
reg [DATAWID-1:0] east15_in151;
reg [DATAWID-1:0] west15_in151;
reg [DATAWID-1:0] north15_in151;
reg [DATAWID-1:0] south15_in151;
reg [DATAWID-1:0] east15_in152;
reg [DATAWID-1:0] west15_in152;
reg [DATAWID-1:0] north15_in152;
reg [DATAWID-1:0] south15_in152;
reg [DATAWID-1:0] east15_in153;
reg [DATAWID-1:0] west15_in153;
reg [DATAWID-1:0] north15_in153;
reg [DATAWID-1:0] south15_in153;
reg [DATAWID-1:0] east15_in154;
reg [DATAWID-1:0] west15_in154;
reg [DATAWID-1:0] north15_in154;
reg [DATAWID-1:0] south15_in154;
reg [DATAWID-1:0] east15_in155;
reg [DATAWID-1:0] west15_in155;
reg [DATAWID-1:0] north15_in155;
reg [DATAWID-1:0] south15_in155;
reg [DATAWID-1:0] east15_in156;
reg [DATAWID-1:0] west15_in156;
reg [DATAWID-1:0] north15_in156;
reg [DATAWID-1:0] south15_in156;
reg [DATAWID-1:0] east15_in157;
reg [DATAWID-1:0] west15_in157;
reg [DATAWID-1:0] north15_in157;
reg [DATAWID-1:0] south15_in157;
reg [DATAWID-1:0] east15_in158;
reg [DATAWID-1:0] west15_in158;
reg [DATAWID-1:0] north15_in158;
reg [DATAWID-1:0] south15_in158;
reg [DATAWID-1:0] east15_in159;
reg [DATAWID-1:0] west15_in159;
reg [DATAWID-1:0] north15_in159;
reg [DATAWID-1:0] south15_in159;
reg [DATAWID-1:0] east15_in1510;
reg [DATAWID-1:0] west15_in1510;
reg [DATAWID-1:0] north15_in1510;
reg [DATAWID-1:0] south15_in1510;
reg [DATAWID-1:0] east15_in1511;
reg [DATAWID-1:0] west15_in1511;
reg [DATAWID-1:0] north15_in1511;
reg [DATAWID-1:0] south15_in1511;
reg [DATAWID-1:0] east15_in1512;
reg [DATAWID-1:0] west15_in1512;
reg [DATAWID-1:0] north15_in1512;
reg [DATAWID-1:0] south15_in1512;
reg [DATAWID-1:0] east15_in1513;
reg [DATAWID-1:0] west15_in1513;
reg [DATAWID-1:0] north15_in1513;
reg [DATAWID-1:0] south15_in1513;
reg [DATAWID-1:0] east15_in1514;
reg [DATAWID-1:0] west15_in1514;
reg [DATAWID-1:0] north15_in1514;
reg [DATAWID-1:0] south15_in1514;
reg [DATAWID-1:0] east15_in1515;
reg [DATAWID-1:0] west15_in1515;
reg [DATAWID-1:0] north15_in1515;
reg [DATAWID-1:0] south15_in1515;
wire [DATAWID-1:0] east0_out00;
wire [DATAWID-1:0] west0_out00;
wire [DATAWID-1:0] north0_out00;
wire [DATAWID-1:0] south0_out00;
wire [DATAWID-1:0] east0_out01;
wire [DATAWID-1:0] west0_out01;
wire [DATAWID-1:0] north0_out01;
wire [DATAWID-1:0] south0_out01;
wire [DATAWID-1:0] east0_out02;
wire [DATAWID-1:0] west0_out02;
wire [DATAWID-1:0] north0_out02;
wire [DATAWID-1:0] south0_out02;
wire [DATAWID-1:0] east0_out03;
wire [DATAWID-1:0] west0_out03;
wire [DATAWID-1:0] north0_out03;
wire [DATAWID-1:0] south0_out03;
wire [DATAWID-1:0] east0_out04;
wire [DATAWID-1:0] west0_out04;
wire [DATAWID-1:0] north0_out04;
wire [DATAWID-1:0] south0_out04;
wire [DATAWID-1:0] east0_out05;
wire [DATAWID-1:0] west0_out05;
wire [DATAWID-1:0] north0_out05;
wire [DATAWID-1:0] south0_out05;
wire [DATAWID-1:0] east0_out06;
wire [DATAWID-1:0] west0_out06;
wire [DATAWID-1:0] north0_out06;
wire [DATAWID-1:0] south0_out06;
wire [DATAWID-1:0] east0_out07;
wire [DATAWID-1:0] west0_out07;
wire [DATAWID-1:0] north0_out07;
wire [DATAWID-1:0] south0_out07;
wire [DATAWID-1:0] east0_out08;
wire [DATAWID-1:0] west0_out08;
wire [DATAWID-1:0] north0_out08;
wire [DATAWID-1:0] south0_out08;
wire [DATAWID-1:0] east0_out09;
wire [DATAWID-1:0] west0_out09;
wire [DATAWID-1:0] north0_out09;
wire [DATAWID-1:0] south0_out09;
wire [DATAWID-1:0] east0_out010;
wire [DATAWID-1:0] west0_out010;
wire [DATAWID-1:0] north0_out010;
wire [DATAWID-1:0] south0_out010;
wire [DATAWID-1:0] east0_out011;
wire [DATAWID-1:0] west0_out011;
wire [DATAWID-1:0] north0_out011;
wire [DATAWID-1:0] south0_out011;
wire [DATAWID-1:0] east0_out012;
wire [DATAWID-1:0] west0_out012;
wire [DATAWID-1:0] north0_out012;
wire [DATAWID-1:0] south0_out012;
wire [DATAWID-1:0] east0_out013;
wire [DATAWID-1:0] west0_out013;
wire [DATAWID-1:0] north0_out013;
wire [DATAWID-1:0] south0_out013;
wire [DATAWID-1:0] east0_out014;
wire [DATAWID-1:0] west0_out014;
wire [DATAWID-1:0] north0_out014;
wire [DATAWID-1:0] south0_out014;
wire [DATAWID-1:0] east0_out015;
wire [DATAWID-1:0] west0_out015;
wire [DATAWID-1:0] north0_out015;
wire [DATAWID-1:0] south0_out015;
wire [DATAWID-1:0] east1_out10;
wire [DATAWID-1:0] west1_out10;
wire [DATAWID-1:0] north1_out10;
wire [DATAWID-1:0] south1_out10;
wire [DATAWID-1:0] east1_out11;
wire [DATAWID-1:0] west1_out11;
wire [DATAWID-1:0] north1_out11;
wire [DATAWID-1:0] south1_out11;
wire [DATAWID-1:0] east1_out12;
wire [DATAWID-1:0] west1_out12;
wire [DATAWID-1:0] north1_out12;
wire [DATAWID-1:0] south1_out12;
wire [DATAWID-1:0] east1_out13;
wire [DATAWID-1:0] west1_out13;
wire [DATAWID-1:0] north1_out13;
wire [DATAWID-1:0] south1_out13;
wire [DATAWID-1:0] east1_out14;
wire [DATAWID-1:0] west1_out14;
wire [DATAWID-1:0] north1_out14;
wire [DATAWID-1:0] south1_out14;
wire [DATAWID-1:0] east1_out15;
wire [DATAWID-1:0] west1_out15;
wire [DATAWID-1:0] north1_out15;
wire [DATAWID-1:0] south1_out15;
wire [DATAWID-1:0] east1_out16;
wire [DATAWID-1:0] west1_out16;
wire [DATAWID-1:0] north1_out16;
wire [DATAWID-1:0] south1_out16;
wire [DATAWID-1:0] east1_out17;
wire [DATAWID-1:0] west1_out17;
wire [DATAWID-1:0] north1_out17;
wire [DATAWID-1:0] south1_out17;
wire [DATAWID-1:0] east1_out18;
wire [DATAWID-1:0] west1_out18;
wire [DATAWID-1:0] north1_out18;
wire [DATAWID-1:0] south1_out18;
wire [DATAWID-1:0] east1_out19;
wire [DATAWID-1:0] west1_out19;
wire [DATAWID-1:0] north1_out19;
wire [DATAWID-1:0] south1_out19;
wire [DATAWID-1:0] east1_out110;
wire [DATAWID-1:0] west1_out110;
wire [DATAWID-1:0] north1_out110;
wire [DATAWID-1:0] south1_out110;
wire [DATAWID-1:0] east1_out111;
wire [DATAWID-1:0] west1_out111;
wire [DATAWID-1:0] north1_out111;
wire [DATAWID-1:0] south1_out111;
wire [DATAWID-1:0] east1_out112;
wire [DATAWID-1:0] west1_out112;
wire [DATAWID-1:0] north1_out112;
wire [DATAWID-1:0] south1_out112;
wire [DATAWID-1:0] east1_out113;
wire [DATAWID-1:0] west1_out113;
wire [DATAWID-1:0] north1_out113;
wire [DATAWID-1:0] south1_out113;
wire [DATAWID-1:0] east1_out114;
wire [DATAWID-1:0] west1_out114;
wire [DATAWID-1:0] north1_out114;
wire [DATAWID-1:0] south1_out114;
wire [DATAWID-1:0] east1_out115;
wire [DATAWID-1:0] west1_out115;
wire [DATAWID-1:0] north1_out115;
wire [DATAWID-1:0] south1_out115;
wire [DATAWID-1:0] east2_out20;
wire [DATAWID-1:0] west2_out20;
wire [DATAWID-1:0] north2_out20;
wire [DATAWID-1:0] south2_out20;
wire [DATAWID-1:0] east2_out21;
wire [DATAWID-1:0] west2_out21;
wire [DATAWID-1:0] north2_out21;
wire [DATAWID-1:0] south2_out21;
wire [DATAWID-1:0] east2_out22;
wire [DATAWID-1:0] west2_out22;
wire [DATAWID-1:0] north2_out22;
wire [DATAWID-1:0] south2_out22;
wire [DATAWID-1:0] east2_out23;
wire [DATAWID-1:0] west2_out23;
wire [DATAWID-1:0] north2_out23;
wire [DATAWID-1:0] south2_out23;
wire [DATAWID-1:0] east2_out24;
wire [DATAWID-1:0] west2_out24;
wire [DATAWID-1:0] north2_out24;
wire [DATAWID-1:0] south2_out24;
wire [DATAWID-1:0] east2_out25;
wire [DATAWID-1:0] west2_out25;
wire [DATAWID-1:0] north2_out25;
wire [DATAWID-1:0] south2_out25;
wire [DATAWID-1:0] east2_out26;
wire [DATAWID-1:0] west2_out26;
wire [DATAWID-1:0] north2_out26;
wire [DATAWID-1:0] south2_out26;
wire [DATAWID-1:0] east2_out27;
wire [DATAWID-1:0] west2_out27;
wire [DATAWID-1:0] north2_out27;
wire [DATAWID-1:0] south2_out27;
wire [DATAWID-1:0] east2_out28;
wire [DATAWID-1:0] west2_out28;
wire [DATAWID-1:0] north2_out28;
wire [DATAWID-1:0] south2_out28;
wire [DATAWID-1:0] east2_out29;
wire [DATAWID-1:0] west2_out29;
wire [DATAWID-1:0] north2_out29;
wire [DATAWID-1:0] south2_out29;
wire [DATAWID-1:0] east2_out210;
wire [DATAWID-1:0] west2_out210;
wire [DATAWID-1:0] north2_out210;
wire [DATAWID-1:0] south2_out210;
wire [DATAWID-1:0] east2_out211;
wire [DATAWID-1:0] west2_out211;
wire [DATAWID-1:0] north2_out211;
wire [DATAWID-1:0] south2_out211;
wire [DATAWID-1:0] east2_out212;
wire [DATAWID-1:0] west2_out212;
wire [DATAWID-1:0] north2_out212;
wire [DATAWID-1:0] south2_out212;
wire [DATAWID-1:0] east2_out213;
wire [DATAWID-1:0] west2_out213;
wire [DATAWID-1:0] north2_out213;
wire [DATAWID-1:0] south2_out213;
wire [DATAWID-1:0] east2_out214;
wire [DATAWID-1:0] west2_out214;
wire [DATAWID-1:0] north2_out214;
wire [DATAWID-1:0] south2_out214;
wire [DATAWID-1:0] east2_out215;
wire [DATAWID-1:0] west2_out215;
wire [DATAWID-1:0] north2_out215;
wire [DATAWID-1:0] south2_out215;
wire [DATAWID-1:0] east3_out30;
wire [DATAWID-1:0] west3_out30;
wire [DATAWID-1:0] north3_out30;
wire [DATAWID-1:0] south3_out30;
wire [DATAWID-1:0] east3_out31;
wire [DATAWID-1:0] west3_out31;
wire [DATAWID-1:0] north3_out31;
wire [DATAWID-1:0] south3_out31;
wire [DATAWID-1:0] east3_out32;
wire [DATAWID-1:0] west3_out32;
wire [DATAWID-1:0] north3_out32;
wire [DATAWID-1:0] south3_out32;
wire [DATAWID-1:0] east3_out33;
wire [DATAWID-1:0] west3_out33;
wire [DATAWID-1:0] north3_out33;
wire [DATAWID-1:0] south3_out33;
wire [DATAWID-1:0] east3_out34;
wire [DATAWID-1:0] west3_out34;
wire [DATAWID-1:0] north3_out34;
wire [DATAWID-1:0] south3_out34;
wire [DATAWID-1:0] east3_out35;
wire [DATAWID-1:0] west3_out35;
wire [DATAWID-1:0] north3_out35;
wire [DATAWID-1:0] south3_out35;
wire [DATAWID-1:0] east3_out36;
wire [DATAWID-1:0] west3_out36;
wire [DATAWID-1:0] north3_out36;
wire [DATAWID-1:0] south3_out36;
wire [DATAWID-1:0] east3_out37;
wire [DATAWID-1:0] west3_out37;
wire [DATAWID-1:0] north3_out37;
wire [DATAWID-1:0] south3_out37;
wire [DATAWID-1:0] east3_out38;
wire [DATAWID-1:0] west3_out38;
wire [DATAWID-1:0] north3_out38;
wire [DATAWID-1:0] south3_out38;
wire [DATAWID-1:0] east3_out39;
wire [DATAWID-1:0] west3_out39;
wire [DATAWID-1:0] north3_out39;
wire [DATAWID-1:0] south3_out39;
wire [DATAWID-1:0] east3_out310;
wire [DATAWID-1:0] west3_out310;
wire [DATAWID-1:0] north3_out310;
wire [DATAWID-1:0] south3_out310;
wire [DATAWID-1:0] east3_out311;
wire [DATAWID-1:0] west3_out311;
wire [DATAWID-1:0] north3_out311;
wire [DATAWID-1:0] south3_out311;
wire [DATAWID-1:0] east3_out312;
wire [DATAWID-1:0] west3_out312;
wire [DATAWID-1:0] north3_out312;
wire [DATAWID-1:0] south3_out312;
wire [DATAWID-1:0] east3_out313;
wire [DATAWID-1:0] west3_out313;
wire [DATAWID-1:0] north3_out313;
wire [DATAWID-1:0] south3_out313;
wire [DATAWID-1:0] east3_out314;
wire [DATAWID-1:0] west3_out314;
wire [DATAWID-1:0] north3_out314;
wire [DATAWID-1:0] south3_out314;
wire [DATAWID-1:0] east3_out315;
wire [DATAWID-1:0] west3_out315;
wire [DATAWID-1:0] north3_out315;
wire [DATAWID-1:0] south3_out315;
wire [DATAWID-1:0] east4_out40;
wire [DATAWID-1:0] west4_out40;
wire [DATAWID-1:0] north4_out40;
wire [DATAWID-1:0] south4_out40;
wire [DATAWID-1:0] east4_out41;
wire [DATAWID-1:0] west4_out41;
wire [DATAWID-1:0] north4_out41;
wire [DATAWID-1:0] south4_out41;
wire [DATAWID-1:0] east4_out42;
wire [DATAWID-1:0] west4_out42;
wire [DATAWID-1:0] north4_out42;
wire [DATAWID-1:0] south4_out42;
wire [DATAWID-1:0] east4_out43;
wire [DATAWID-1:0] west4_out43;
wire [DATAWID-1:0] north4_out43;
wire [DATAWID-1:0] south4_out43;
wire [DATAWID-1:0] east4_out44;
wire [DATAWID-1:0] west4_out44;
wire [DATAWID-1:0] north4_out44;
wire [DATAWID-1:0] south4_out44;
wire [DATAWID-1:0] east4_out45;
wire [DATAWID-1:0] west4_out45;
wire [DATAWID-1:0] north4_out45;
wire [DATAWID-1:0] south4_out45;
wire [DATAWID-1:0] east4_out46;
wire [DATAWID-1:0] west4_out46;
wire [DATAWID-1:0] north4_out46;
wire [DATAWID-1:0] south4_out46;
wire [DATAWID-1:0] east4_out47;
wire [DATAWID-1:0] west4_out47;
wire [DATAWID-1:0] north4_out47;
wire [DATAWID-1:0] south4_out47;
wire [DATAWID-1:0] east4_out48;
wire [DATAWID-1:0] west4_out48;
wire [DATAWID-1:0] north4_out48;
wire [DATAWID-1:0] south4_out48;
wire [DATAWID-1:0] east4_out49;
wire [DATAWID-1:0] west4_out49;
wire [DATAWID-1:0] north4_out49;
wire [DATAWID-1:0] south4_out49;
wire [DATAWID-1:0] east4_out410;
wire [DATAWID-1:0] west4_out410;
wire [DATAWID-1:0] north4_out410;
wire [DATAWID-1:0] south4_out410;
wire [DATAWID-1:0] east4_out411;
wire [DATAWID-1:0] west4_out411;
wire [DATAWID-1:0] north4_out411;
wire [DATAWID-1:0] south4_out411;
wire [DATAWID-1:0] east4_out412;
wire [DATAWID-1:0] west4_out412;
wire [DATAWID-1:0] north4_out412;
wire [DATAWID-1:0] south4_out412;
wire [DATAWID-1:0] east4_out413;
wire [DATAWID-1:0] west4_out413;
wire [DATAWID-1:0] north4_out413;
wire [DATAWID-1:0] south4_out413;
wire [DATAWID-1:0] east4_out414;
wire [DATAWID-1:0] west4_out414;
wire [DATAWID-1:0] north4_out414;
wire [DATAWID-1:0] south4_out414;
wire [DATAWID-1:0] east4_out415;
wire [DATAWID-1:0] west4_out415;
wire [DATAWID-1:0] north4_out415;
wire [DATAWID-1:0] south4_out415;
wire [DATAWID-1:0] east5_out50;
wire [DATAWID-1:0] west5_out50;
wire [DATAWID-1:0] north5_out50;
wire [DATAWID-1:0] south5_out50;
wire [DATAWID-1:0] east5_out51;
wire [DATAWID-1:0] west5_out51;
wire [DATAWID-1:0] north5_out51;
wire [DATAWID-1:0] south5_out51;
wire [DATAWID-1:0] east5_out52;
wire [DATAWID-1:0] west5_out52;
wire [DATAWID-1:0] north5_out52;
wire [DATAWID-1:0] south5_out52;
wire [DATAWID-1:0] east5_out53;
wire [DATAWID-1:0] west5_out53;
wire [DATAWID-1:0] north5_out53;
wire [DATAWID-1:0] south5_out53;
wire [DATAWID-1:0] east5_out54;
wire [DATAWID-1:0] west5_out54;
wire [DATAWID-1:0] north5_out54;
wire [DATAWID-1:0] south5_out54;
wire [DATAWID-1:0] east5_out55;
wire [DATAWID-1:0] west5_out55;
wire [DATAWID-1:0] north5_out55;
wire [DATAWID-1:0] south5_out55;
wire [DATAWID-1:0] east5_out56;
wire [DATAWID-1:0] west5_out56;
wire [DATAWID-1:0] north5_out56;
wire [DATAWID-1:0] south5_out56;
wire [DATAWID-1:0] east5_out57;
wire [DATAWID-1:0] west5_out57;
wire [DATAWID-1:0] north5_out57;
wire [DATAWID-1:0] south5_out57;
wire [DATAWID-1:0] east5_out58;
wire [DATAWID-1:0] west5_out58;
wire [DATAWID-1:0] north5_out58;
wire [DATAWID-1:0] south5_out58;
wire [DATAWID-1:0] east5_out59;
wire [DATAWID-1:0] west5_out59;
wire [DATAWID-1:0] north5_out59;
wire [DATAWID-1:0] south5_out59;
wire [DATAWID-1:0] east5_out510;
wire [DATAWID-1:0] west5_out510;
wire [DATAWID-1:0] north5_out510;
wire [DATAWID-1:0] south5_out510;
wire [DATAWID-1:0] east5_out511;
wire [DATAWID-1:0] west5_out511;
wire [DATAWID-1:0] north5_out511;
wire [DATAWID-1:0] south5_out511;
wire [DATAWID-1:0] east5_out512;
wire [DATAWID-1:0] west5_out512;
wire [DATAWID-1:0] north5_out512;
wire [DATAWID-1:0] south5_out512;
wire [DATAWID-1:0] east5_out513;
wire [DATAWID-1:0] west5_out513;
wire [DATAWID-1:0] north5_out513;
wire [DATAWID-1:0] south5_out513;
wire [DATAWID-1:0] east5_out514;
wire [DATAWID-1:0] west5_out514;
wire [DATAWID-1:0] north5_out514;
wire [DATAWID-1:0] south5_out514;
wire [DATAWID-1:0] east5_out515;
wire [DATAWID-1:0] west5_out515;
wire [DATAWID-1:0] north5_out515;
wire [DATAWID-1:0] south5_out515;
wire [DATAWID-1:0] east6_out60;
wire [DATAWID-1:0] west6_out60;
wire [DATAWID-1:0] north6_out60;
wire [DATAWID-1:0] south6_out60;
wire [DATAWID-1:0] east6_out61;
wire [DATAWID-1:0] west6_out61;
wire [DATAWID-1:0] north6_out61;
wire [DATAWID-1:0] south6_out61;
wire [DATAWID-1:0] east6_out62;
wire [DATAWID-1:0] west6_out62;
wire [DATAWID-1:0] north6_out62;
wire [DATAWID-1:0] south6_out62;
wire [DATAWID-1:0] east6_out63;
wire [DATAWID-1:0] west6_out63;
wire [DATAWID-1:0] north6_out63;
wire [DATAWID-1:0] south6_out63;
wire [DATAWID-1:0] east6_out64;
wire [DATAWID-1:0] west6_out64;
wire [DATAWID-1:0] north6_out64;
wire [DATAWID-1:0] south6_out64;
wire [DATAWID-1:0] east6_out65;
wire [DATAWID-1:0] west6_out65;
wire [DATAWID-1:0] north6_out65;
wire [DATAWID-1:0] south6_out65;
wire [DATAWID-1:0] east6_out66;
wire [DATAWID-1:0] west6_out66;
wire [DATAWID-1:0] north6_out66;
wire [DATAWID-1:0] south6_out66;
wire [DATAWID-1:0] east6_out67;
wire [DATAWID-1:0] west6_out67;
wire [DATAWID-1:0] north6_out67;
wire [DATAWID-1:0] south6_out67;
wire [DATAWID-1:0] east6_out68;
wire [DATAWID-1:0] west6_out68;
wire [DATAWID-1:0] north6_out68;
wire [DATAWID-1:0] south6_out68;
wire [DATAWID-1:0] east6_out69;
wire [DATAWID-1:0] west6_out69;
wire [DATAWID-1:0] north6_out69;
wire [DATAWID-1:0] south6_out69;
wire [DATAWID-1:0] east6_out610;
wire [DATAWID-1:0] west6_out610;
wire [DATAWID-1:0] north6_out610;
wire [DATAWID-1:0] south6_out610;
wire [DATAWID-1:0] east6_out611;
wire [DATAWID-1:0] west6_out611;
wire [DATAWID-1:0] north6_out611;
wire [DATAWID-1:0] south6_out611;
wire [DATAWID-1:0] east6_out612;
wire [DATAWID-1:0] west6_out612;
wire [DATAWID-1:0] north6_out612;
wire [DATAWID-1:0] south6_out612;
wire [DATAWID-1:0] east6_out613;
wire [DATAWID-1:0] west6_out613;
wire [DATAWID-1:0] north6_out613;
wire [DATAWID-1:0] south6_out613;
wire [DATAWID-1:0] east6_out614;
wire [DATAWID-1:0] west6_out614;
wire [DATAWID-1:0] north6_out614;
wire [DATAWID-1:0] south6_out614;
wire [DATAWID-1:0] east6_out615;
wire [DATAWID-1:0] west6_out615;
wire [DATAWID-1:0] north6_out615;
wire [DATAWID-1:0] south6_out615;
wire [DATAWID-1:0] east7_out70;
wire [DATAWID-1:0] west7_out70;
wire [DATAWID-1:0] north7_out70;
wire [DATAWID-1:0] south7_out70;
wire [DATAWID-1:0] east7_out71;
wire [DATAWID-1:0] west7_out71;
wire [DATAWID-1:0] north7_out71;
wire [DATAWID-1:0] south7_out71;
wire [DATAWID-1:0] east7_out72;
wire [DATAWID-1:0] west7_out72;
wire [DATAWID-1:0] north7_out72;
wire [DATAWID-1:0] south7_out72;
wire [DATAWID-1:0] east7_out73;
wire [DATAWID-1:0] west7_out73;
wire [DATAWID-1:0] north7_out73;
wire [DATAWID-1:0] south7_out73;
wire [DATAWID-1:0] east7_out74;
wire [DATAWID-1:0] west7_out74;
wire [DATAWID-1:0] north7_out74;
wire [DATAWID-1:0] south7_out74;
wire [DATAWID-1:0] east7_out75;
wire [DATAWID-1:0] west7_out75;
wire [DATAWID-1:0] north7_out75;
wire [DATAWID-1:0] south7_out75;
wire [DATAWID-1:0] east7_out76;
wire [DATAWID-1:0] west7_out76;
wire [DATAWID-1:0] north7_out76;
wire [DATAWID-1:0] south7_out76;
wire [DATAWID-1:0] east7_out77;
wire [DATAWID-1:0] west7_out77;
wire [DATAWID-1:0] north7_out77;
wire [DATAWID-1:0] south7_out77;
wire [DATAWID-1:0] east7_out78;
wire [DATAWID-1:0] west7_out78;
wire [DATAWID-1:0] north7_out78;
wire [DATAWID-1:0] south7_out78;
wire [DATAWID-1:0] east7_out79;
wire [DATAWID-1:0] west7_out79;
wire [DATAWID-1:0] north7_out79;
wire [DATAWID-1:0] south7_out79;
wire [DATAWID-1:0] east7_out710;
wire [DATAWID-1:0] west7_out710;
wire [DATAWID-1:0] north7_out710;
wire [DATAWID-1:0] south7_out710;
wire [DATAWID-1:0] east7_out711;
wire [DATAWID-1:0] west7_out711;
wire [DATAWID-1:0] north7_out711;
wire [DATAWID-1:0] south7_out711;
wire [DATAWID-1:0] east7_out712;
wire [DATAWID-1:0] west7_out712;
wire [DATAWID-1:0] north7_out712;
wire [DATAWID-1:0] south7_out712;
wire [DATAWID-1:0] east7_out713;
wire [DATAWID-1:0] west7_out713;
wire [DATAWID-1:0] north7_out713;
wire [DATAWID-1:0] south7_out713;
wire [DATAWID-1:0] east7_out714;
wire [DATAWID-1:0] west7_out714;
wire [DATAWID-1:0] north7_out714;
wire [DATAWID-1:0] south7_out714;
wire [DATAWID-1:0] east7_out715;
wire [DATAWID-1:0] west7_out715;
wire [DATAWID-1:0] north7_out715;
wire [DATAWID-1:0] south7_out715;
wire [DATAWID-1:0] east8_out80;
wire [DATAWID-1:0] west8_out80;
wire [DATAWID-1:0] north8_out80;
wire [DATAWID-1:0] south8_out80;
wire [DATAWID-1:0] east8_out81;
wire [DATAWID-1:0] west8_out81;
wire [DATAWID-1:0] north8_out81;
wire [DATAWID-1:0] south8_out81;
wire [DATAWID-1:0] east8_out82;
wire [DATAWID-1:0] west8_out82;
wire [DATAWID-1:0] north8_out82;
wire [DATAWID-1:0] south8_out82;
wire [DATAWID-1:0] east8_out83;
wire [DATAWID-1:0] west8_out83;
wire [DATAWID-1:0] north8_out83;
wire [DATAWID-1:0] south8_out83;
wire [DATAWID-1:0] east8_out84;
wire [DATAWID-1:0] west8_out84;
wire [DATAWID-1:0] north8_out84;
wire [DATAWID-1:0] south8_out84;
wire [DATAWID-1:0] east8_out85;
wire [DATAWID-1:0] west8_out85;
wire [DATAWID-1:0] north8_out85;
wire [DATAWID-1:0] south8_out85;
wire [DATAWID-1:0] east8_out86;
wire [DATAWID-1:0] west8_out86;
wire [DATAWID-1:0] north8_out86;
wire [DATAWID-1:0] south8_out86;
wire [DATAWID-1:0] east8_out87;
wire [DATAWID-1:0] west8_out87;
wire [DATAWID-1:0] north8_out87;
wire [DATAWID-1:0] south8_out87;
wire [DATAWID-1:0] east8_out88;
wire [DATAWID-1:0] west8_out88;
wire [DATAWID-1:0] north8_out88;
wire [DATAWID-1:0] south8_out88;
wire [DATAWID-1:0] east8_out89;
wire [DATAWID-1:0] west8_out89;
wire [DATAWID-1:0] north8_out89;
wire [DATAWID-1:0] south8_out89;
wire [DATAWID-1:0] east8_out810;
wire [DATAWID-1:0] west8_out810;
wire [DATAWID-1:0] north8_out810;
wire [DATAWID-1:0] south8_out810;
wire [DATAWID-1:0] east8_out811;
wire [DATAWID-1:0] west8_out811;
wire [DATAWID-1:0] north8_out811;
wire [DATAWID-1:0] south8_out811;
wire [DATAWID-1:0] east8_out812;
wire [DATAWID-1:0] west8_out812;
wire [DATAWID-1:0] north8_out812;
wire [DATAWID-1:0] south8_out812;
wire [DATAWID-1:0] east8_out813;
wire [DATAWID-1:0] west8_out813;
wire [DATAWID-1:0] north8_out813;
wire [DATAWID-1:0] south8_out813;
wire [DATAWID-1:0] east8_out814;
wire [DATAWID-1:0] west8_out814;
wire [DATAWID-1:0] north8_out814;
wire [DATAWID-1:0] south8_out814;
wire [DATAWID-1:0] east8_out815;
wire [DATAWID-1:0] west8_out815;
wire [DATAWID-1:0] north8_out815;
wire [DATAWID-1:0] south8_out815;
wire [DATAWID-1:0] east9_out90;
wire [DATAWID-1:0] west9_out90;
wire [DATAWID-1:0] north9_out90;
wire [DATAWID-1:0] south9_out90;
wire [DATAWID-1:0] east9_out91;
wire [DATAWID-1:0] west9_out91;
wire [DATAWID-1:0] north9_out91;
wire [DATAWID-1:0] south9_out91;
wire [DATAWID-1:0] east9_out92;
wire [DATAWID-1:0] west9_out92;
wire [DATAWID-1:0] north9_out92;
wire [DATAWID-1:0] south9_out92;
wire [DATAWID-1:0] east9_out93;
wire [DATAWID-1:0] west9_out93;
wire [DATAWID-1:0] north9_out93;
wire [DATAWID-1:0] south9_out93;
wire [DATAWID-1:0] east9_out94;
wire [DATAWID-1:0] west9_out94;
wire [DATAWID-1:0] north9_out94;
wire [DATAWID-1:0] south9_out94;
wire [DATAWID-1:0] east9_out95;
wire [DATAWID-1:0] west9_out95;
wire [DATAWID-1:0] north9_out95;
wire [DATAWID-1:0] south9_out95;
wire [DATAWID-1:0] east9_out96;
wire [DATAWID-1:0] west9_out96;
wire [DATAWID-1:0] north9_out96;
wire [DATAWID-1:0] south9_out96;
wire [DATAWID-1:0] east9_out97;
wire [DATAWID-1:0] west9_out97;
wire [DATAWID-1:0] north9_out97;
wire [DATAWID-1:0] south9_out97;
wire [DATAWID-1:0] east9_out98;
wire [DATAWID-1:0] west9_out98;
wire [DATAWID-1:0] north9_out98;
wire [DATAWID-1:0] south9_out98;
wire [DATAWID-1:0] east9_out99;
wire [DATAWID-1:0] west9_out99;
wire [DATAWID-1:0] north9_out99;
wire [DATAWID-1:0] south9_out99;
wire [DATAWID-1:0] east9_out910;
wire [DATAWID-1:0] west9_out910;
wire [DATAWID-1:0] north9_out910;
wire [DATAWID-1:0] south9_out910;
wire [DATAWID-1:0] east9_out911;
wire [DATAWID-1:0] west9_out911;
wire [DATAWID-1:0] north9_out911;
wire [DATAWID-1:0] south9_out911;
wire [DATAWID-1:0] east9_out912;
wire [DATAWID-1:0] west9_out912;
wire [DATAWID-1:0] north9_out912;
wire [DATAWID-1:0] south9_out912;
wire [DATAWID-1:0] east9_out913;
wire [DATAWID-1:0] west9_out913;
wire [DATAWID-1:0] north9_out913;
wire [DATAWID-1:0] south9_out913;
wire [DATAWID-1:0] east9_out914;
wire [DATAWID-1:0] west9_out914;
wire [DATAWID-1:0] north9_out914;
wire [DATAWID-1:0] south9_out914;
wire [DATAWID-1:0] east9_out915;
wire [DATAWID-1:0] west9_out915;
wire [DATAWID-1:0] north9_out915;
wire [DATAWID-1:0] south9_out915;
wire [DATAWID-1:0] east10_out100;
wire [DATAWID-1:0] west10_out100;
wire [DATAWID-1:0] north10_out100;
wire [DATAWID-1:0] south10_out100;
wire [DATAWID-1:0] east10_out101;
wire [DATAWID-1:0] west10_out101;
wire [DATAWID-1:0] north10_out101;
wire [DATAWID-1:0] south10_out101;
wire [DATAWID-1:0] east10_out102;
wire [DATAWID-1:0] west10_out102;
wire [DATAWID-1:0] north10_out102;
wire [DATAWID-1:0] south10_out102;
wire [DATAWID-1:0] east10_out103;
wire [DATAWID-1:0] west10_out103;
wire [DATAWID-1:0] north10_out103;
wire [DATAWID-1:0] south10_out103;
wire [DATAWID-1:0] east10_out104;
wire [DATAWID-1:0] west10_out104;
wire [DATAWID-1:0] north10_out104;
wire [DATAWID-1:0] south10_out104;
wire [DATAWID-1:0] east10_out105;
wire [DATAWID-1:0] west10_out105;
wire [DATAWID-1:0] north10_out105;
wire [DATAWID-1:0] south10_out105;
wire [DATAWID-1:0] east10_out106;
wire [DATAWID-1:0] west10_out106;
wire [DATAWID-1:0] north10_out106;
wire [DATAWID-1:0] south10_out106;
wire [DATAWID-1:0] east10_out107;
wire [DATAWID-1:0] west10_out107;
wire [DATAWID-1:0] north10_out107;
wire [DATAWID-1:0] south10_out107;
wire [DATAWID-1:0] east10_out108;
wire [DATAWID-1:0] west10_out108;
wire [DATAWID-1:0] north10_out108;
wire [DATAWID-1:0] south10_out108;
wire [DATAWID-1:0] east10_out109;
wire [DATAWID-1:0] west10_out109;
wire [DATAWID-1:0] north10_out109;
wire [DATAWID-1:0] south10_out109;
wire [DATAWID-1:0] east10_out1010;
wire [DATAWID-1:0] west10_out1010;
wire [DATAWID-1:0] north10_out1010;
wire [DATAWID-1:0] south10_out1010;
wire [DATAWID-1:0] east10_out1011;
wire [DATAWID-1:0] west10_out1011;
wire [DATAWID-1:0] north10_out1011;
wire [DATAWID-1:0] south10_out1011;
wire [DATAWID-1:0] east10_out1012;
wire [DATAWID-1:0] west10_out1012;
wire [DATAWID-1:0] north10_out1012;
wire [DATAWID-1:0] south10_out1012;
wire [DATAWID-1:0] east10_out1013;
wire [DATAWID-1:0] west10_out1013;
wire [DATAWID-1:0] north10_out1013;
wire [DATAWID-1:0] south10_out1013;
wire [DATAWID-1:0] east10_out1014;
wire [DATAWID-1:0] west10_out1014;
wire [DATAWID-1:0] north10_out1014;
wire [DATAWID-1:0] south10_out1014;
wire [DATAWID-1:0] east10_out1015;
wire [DATAWID-1:0] west10_out1015;
wire [DATAWID-1:0] north10_out1015;
wire [DATAWID-1:0] south10_out1015;
wire [DATAWID-1:0] east11_out110;
wire [DATAWID-1:0] west11_out110;
wire [DATAWID-1:0] north11_out110;
wire [DATAWID-1:0] south11_out110;
wire [DATAWID-1:0] east11_out111;
wire [DATAWID-1:0] west11_out111;
wire [DATAWID-1:0] north11_out111;
wire [DATAWID-1:0] south11_out111;
wire [DATAWID-1:0] east11_out112;
wire [DATAWID-1:0] west11_out112;
wire [DATAWID-1:0] north11_out112;
wire [DATAWID-1:0] south11_out112;
wire [DATAWID-1:0] east11_out113;
wire [DATAWID-1:0] west11_out113;
wire [DATAWID-1:0] north11_out113;
wire [DATAWID-1:0] south11_out113;
wire [DATAWID-1:0] east11_out114;
wire [DATAWID-1:0] west11_out114;
wire [DATAWID-1:0] north11_out114;
wire [DATAWID-1:0] south11_out114;
wire [DATAWID-1:0] east11_out115;
wire [DATAWID-1:0] west11_out115;
wire [DATAWID-1:0] north11_out115;
wire [DATAWID-1:0] south11_out115;
wire [DATAWID-1:0] east11_out116;
wire [DATAWID-1:0] west11_out116;
wire [DATAWID-1:0] north11_out116;
wire [DATAWID-1:0] south11_out116;
wire [DATAWID-1:0] east11_out117;
wire [DATAWID-1:0] west11_out117;
wire [DATAWID-1:0] north11_out117;
wire [DATAWID-1:0] south11_out117;
wire [DATAWID-1:0] east11_out118;
wire [DATAWID-1:0] west11_out118;
wire [DATAWID-1:0] north11_out118;
wire [DATAWID-1:0] south11_out118;
wire [DATAWID-1:0] east11_out119;
wire [DATAWID-1:0] west11_out119;
wire [DATAWID-1:0] north11_out119;
wire [DATAWID-1:0] south11_out119;
wire [DATAWID-1:0] east11_out1110;
wire [DATAWID-1:0] west11_out1110;
wire [DATAWID-1:0] north11_out1110;
wire [DATAWID-1:0] south11_out1110;
wire [DATAWID-1:0] east11_out1111;
wire [DATAWID-1:0] west11_out1111;
wire [DATAWID-1:0] north11_out1111;
wire [DATAWID-1:0] south11_out1111;
wire [DATAWID-1:0] east11_out1112;
wire [DATAWID-1:0] west11_out1112;
wire [DATAWID-1:0] north11_out1112;
wire [DATAWID-1:0] south11_out1112;
wire [DATAWID-1:0] east11_out1113;
wire [DATAWID-1:0] west11_out1113;
wire [DATAWID-1:0] north11_out1113;
wire [DATAWID-1:0] south11_out1113;
wire [DATAWID-1:0] east11_out1114;
wire [DATAWID-1:0] west11_out1114;
wire [DATAWID-1:0] north11_out1114;
wire [DATAWID-1:0] south11_out1114;
wire [DATAWID-1:0] east11_out1115;
wire [DATAWID-1:0] west11_out1115;
wire [DATAWID-1:0] north11_out1115;
wire [DATAWID-1:0] south11_out1115;
wire [DATAWID-1:0] east12_out120;
wire [DATAWID-1:0] west12_out120;
wire [DATAWID-1:0] north12_out120;
wire [DATAWID-1:0] south12_out120;
wire [DATAWID-1:0] east12_out121;
wire [DATAWID-1:0] west12_out121;
wire [DATAWID-1:0] north12_out121;
wire [DATAWID-1:0] south12_out121;
wire [DATAWID-1:0] east12_out122;
wire [DATAWID-1:0] west12_out122;
wire [DATAWID-1:0] north12_out122;
wire [DATAWID-1:0] south12_out122;
wire [DATAWID-1:0] east12_out123;
wire [DATAWID-1:0] west12_out123;
wire [DATAWID-1:0] north12_out123;
wire [DATAWID-1:0] south12_out123;
wire [DATAWID-1:0] east12_out124;
wire [DATAWID-1:0] west12_out124;
wire [DATAWID-1:0] north12_out124;
wire [DATAWID-1:0] south12_out124;
wire [DATAWID-1:0] east12_out125;
wire [DATAWID-1:0] west12_out125;
wire [DATAWID-1:0] north12_out125;
wire [DATAWID-1:0] south12_out125;
wire [DATAWID-1:0] east12_out126;
wire [DATAWID-1:0] west12_out126;
wire [DATAWID-1:0] north12_out126;
wire [DATAWID-1:0] south12_out126;
wire [DATAWID-1:0] east12_out127;
wire [DATAWID-1:0] west12_out127;
wire [DATAWID-1:0] north12_out127;
wire [DATAWID-1:0] south12_out127;
wire [DATAWID-1:0] east12_out128;
wire [DATAWID-1:0] west12_out128;
wire [DATAWID-1:0] north12_out128;
wire [DATAWID-1:0] south12_out128;
wire [DATAWID-1:0] east12_out129;
wire [DATAWID-1:0] west12_out129;
wire [DATAWID-1:0] north12_out129;
wire [DATAWID-1:0] south12_out129;
wire [DATAWID-1:0] east12_out1210;
wire [DATAWID-1:0] west12_out1210;
wire [DATAWID-1:0] north12_out1210;
wire [DATAWID-1:0] south12_out1210;
wire [DATAWID-1:0] east12_out1211;
wire [DATAWID-1:0] west12_out1211;
wire [DATAWID-1:0] north12_out1211;
wire [DATAWID-1:0] south12_out1211;
wire [DATAWID-1:0] east12_out1212;
wire [DATAWID-1:0] west12_out1212;
wire [DATAWID-1:0] north12_out1212;
wire [DATAWID-1:0] south12_out1212;
wire [DATAWID-1:0] east12_out1213;
wire [DATAWID-1:0] west12_out1213;
wire [DATAWID-1:0] north12_out1213;
wire [DATAWID-1:0] south12_out1213;
wire [DATAWID-1:0] east12_out1214;
wire [DATAWID-1:0] west12_out1214;
wire [DATAWID-1:0] north12_out1214;
wire [DATAWID-1:0] south12_out1214;
wire [DATAWID-1:0] east12_out1215;
wire [DATAWID-1:0] west12_out1215;
wire [DATAWID-1:0] north12_out1215;
wire [DATAWID-1:0] south12_out1215;
wire [DATAWID-1:0] east13_out130;
wire [DATAWID-1:0] west13_out130;
wire [DATAWID-1:0] north13_out130;
wire [DATAWID-1:0] south13_out130;
wire [DATAWID-1:0] east13_out131;
wire [DATAWID-1:0] west13_out131;
wire [DATAWID-1:0] north13_out131;
wire [DATAWID-1:0] south13_out131;
wire [DATAWID-1:0] east13_out132;
wire [DATAWID-1:0] west13_out132;
wire [DATAWID-1:0] north13_out132;
wire [DATAWID-1:0] south13_out132;
wire [DATAWID-1:0] east13_out133;
wire [DATAWID-1:0] west13_out133;
wire [DATAWID-1:0] north13_out133;
wire [DATAWID-1:0] south13_out133;
wire [DATAWID-1:0] east13_out134;
wire [DATAWID-1:0] west13_out134;
wire [DATAWID-1:0] north13_out134;
wire [DATAWID-1:0] south13_out134;
wire [DATAWID-1:0] east13_out135;
wire [DATAWID-1:0] west13_out135;
wire [DATAWID-1:0] north13_out135;
wire [DATAWID-1:0] south13_out135;
wire [DATAWID-1:0] east13_out136;
wire [DATAWID-1:0] west13_out136;
wire [DATAWID-1:0] north13_out136;
wire [DATAWID-1:0] south13_out136;
wire [DATAWID-1:0] east13_out137;
wire [DATAWID-1:0] west13_out137;
wire [DATAWID-1:0] north13_out137;
wire [DATAWID-1:0] south13_out137;
wire [DATAWID-1:0] east13_out138;
wire [DATAWID-1:0] west13_out138;
wire [DATAWID-1:0] north13_out138;
wire [DATAWID-1:0] south13_out138;
wire [DATAWID-1:0] east13_out139;
wire [DATAWID-1:0] west13_out139;
wire [DATAWID-1:0] north13_out139;
wire [DATAWID-1:0] south13_out139;
wire [DATAWID-1:0] east13_out1310;
wire [DATAWID-1:0] west13_out1310;
wire [DATAWID-1:0] north13_out1310;
wire [DATAWID-1:0] south13_out1310;
wire [DATAWID-1:0] east13_out1311;
wire [DATAWID-1:0] west13_out1311;
wire [DATAWID-1:0] north13_out1311;
wire [DATAWID-1:0] south13_out1311;
wire [DATAWID-1:0] east13_out1312;
wire [DATAWID-1:0] west13_out1312;
wire [DATAWID-1:0] north13_out1312;
wire [DATAWID-1:0] south13_out1312;
wire [DATAWID-1:0] east13_out1313;
wire [DATAWID-1:0] west13_out1313;
wire [DATAWID-1:0] north13_out1313;
wire [DATAWID-1:0] south13_out1313;
wire [DATAWID-1:0] east13_out1314;
wire [DATAWID-1:0] west13_out1314;
wire [DATAWID-1:0] north13_out1314;
wire [DATAWID-1:0] south13_out1314;
wire [DATAWID-1:0] east13_out1315;
wire [DATAWID-1:0] west13_out1315;
wire [DATAWID-1:0] north13_out1315;
wire [DATAWID-1:0] south13_out1315;
wire [DATAWID-1:0] east14_out140;
wire [DATAWID-1:0] west14_out140;
wire [DATAWID-1:0] north14_out140;
wire [DATAWID-1:0] south14_out140;
wire [DATAWID-1:0] east14_out141;
wire [DATAWID-1:0] west14_out141;
wire [DATAWID-1:0] north14_out141;
wire [DATAWID-1:0] south14_out141;
wire [DATAWID-1:0] east14_out142;
wire [DATAWID-1:0] west14_out142;
wire [DATAWID-1:0] north14_out142;
wire [DATAWID-1:0] south14_out142;
wire [DATAWID-1:0] east14_out143;
wire [DATAWID-1:0] west14_out143;
wire [DATAWID-1:0] north14_out143;
wire [DATAWID-1:0] south14_out143;
wire [DATAWID-1:0] east14_out144;
wire [DATAWID-1:0] west14_out144;
wire [DATAWID-1:0] north14_out144;
wire [DATAWID-1:0] south14_out144;
wire [DATAWID-1:0] east14_out145;
wire [DATAWID-1:0] west14_out145;
wire [DATAWID-1:0] north14_out145;
wire [DATAWID-1:0] south14_out145;
wire [DATAWID-1:0] east14_out146;
wire [DATAWID-1:0] west14_out146;
wire [DATAWID-1:0] north14_out146;
wire [DATAWID-1:0] south14_out146;
wire [DATAWID-1:0] east14_out147;
wire [DATAWID-1:0] west14_out147;
wire [DATAWID-1:0] north14_out147;
wire [DATAWID-1:0] south14_out147;
wire [DATAWID-1:0] east14_out148;
wire [DATAWID-1:0] west14_out148;
wire [DATAWID-1:0] north14_out148;
wire [DATAWID-1:0] south14_out148;
wire [DATAWID-1:0] east14_out149;
wire [DATAWID-1:0] west14_out149;
wire [DATAWID-1:0] north14_out149;
wire [DATAWID-1:0] south14_out149;
wire [DATAWID-1:0] east14_out1410;
wire [DATAWID-1:0] west14_out1410;
wire [DATAWID-1:0] north14_out1410;
wire [DATAWID-1:0] south14_out1410;
wire [DATAWID-1:0] east14_out1411;
wire [DATAWID-1:0] west14_out1411;
wire [DATAWID-1:0] north14_out1411;
wire [DATAWID-1:0] south14_out1411;
wire [DATAWID-1:0] east14_out1412;
wire [DATAWID-1:0] west14_out1412;
wire [DATAWID-1:0] north14_out1412;
wire [DATAWID-1:0] south14_out1412;
wire [DATAWID-1:0] east14_out1413;
wire [DATAWID-1:0] west14_out1413;
wire [DATAWID-1:0] north14_out1413;
wire [DATAWID-1:0] south14_out1413;
wire [DATAWID-1:0] east14_out1414;
wire [DATAWID-1:0] west14_out1414;
wire [DATAWID-1:0] north14_out1414;
wire [DATAWID-1:0] south14_out1414;
wire [DATAWID-1:0] east14_out1415;
wire [DATAWID-1:0] west14_out1415;
wire [DATAWID-1:0] north14_out1415;
wire [DATAWID-1:0] south14_out1415;
wire [DATAWID-1:0] east15_out150;
wire [DATAWID-1:0] west15_out150;
wire [DATAWID-1:0] north15_out150;
wire [DATAWID-1:0] south15_out150;
wire [DATAWID-1:0] east15_out151;
wire [DATAWID-1:0] west15_out151;
wire [DATAWID-1:0] north15_out151;
wire [DATAWID-1:0] south15_out151;
wire [DATAWID-1:0] east15_out152;
wire [DATAWID-1:0] west15_out152;
wire [DATAWID-1:0] north15_out152;
wire [DATAWID-1:0] south15_out152;
wire [DATAWID-1:0] east15_out153;
wire [DATAWID-1:0] west15_out153;
wire [DATAWID-1:0] north15_out153;
wire [DATAWID-1:0] south15_out153;
wire [DATAWID-1:0] east15_out154;
wire [DATAWID-1:0] west15_out154;
wire [DATAWID-1:0] north15_out154;
wire [DATAWID-1:0] south15_out154;
wire [DATAWID-1:0] east15_out155;
wire [DATAWID-1:0] west15_out155;
wire [DATAWID-1:0] north15_out155;
wire [DATAWID-1:0] south15_out155;
wire [DATAWID-1:0] east15_out156;
wire [DATAWID-1:0] west15_out156;
wire [DATAWID-1:0] north15_out156;
wire [DATAWID-1:0] south15_out156;
wire [DATAWID-1:0] east15_out157;
wire [DATAWID-1:0] west15_out157;
wire [DATAWID-1:0] north15_out157;
wire [DATAWID-1:0] south15_out157;
wire [DATAWID-1:0] east15_out158;
wire [DATAWID-1:0] west15_out158;
wire [DATAWID-1:0] north15_out158;
wire [DATAWID-1:0] south15_out158;
wire [DATAWID-1:0] east15_out159;
wire [DATAWID-1:0] west15_out159;
wire [DATAWID-1:0] north15_out159;
wire [DATAWID-1:0] south15_out159;
wire [DATAWID-1:0] east15_out1510;
wire [DATAWID-1:0] west15_out1510;
wire [DATAWID-1:0] north15_out1510;
wire [DATAWID-1:0] south15_out1510;
wire [DATAWID-1:0] east15_out1511;
wire [DATAWID-1:0] west15_out1511;
wire [DATAWID-1:0] north15_out1511;
wire [DATAWID-1:0] south15_out1511;
wire [DATAWID-1:0] east15_out1512;
wire [DATAWID-1:0] west15_out1512;
wire [DATAWID-1:0] north15_out1512;
wire [DATAWID-1:0] south15_out1512;
wire [DATAWID-1:0] east15_out1513;
wire [DATAWID-1:0] west15_out1513;
wire [DATAWID-1:0] north15_out1513;
wire [DATAWID-1:0] south15_out1513;
wire [DATAWID-1:0] east15_out1514;
wire [DATAWID-1:0] west15_out1514;
wire [DATAWID-1:0] north15_out1514;
wire [DATAWID-1:0] south15_out1514;
wire [DATAWID-1:0] east15_out1515;
wire [DATAWID-1:0] west15_out1515;
wire [DATAWID-1:0] north15_out1515;
wire [DATAWID-1:0] south15_out1515;
router r000
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in00),
.i01(east0_in00),
.i02(west0_in00),
.i03(north0_in00),
.i04(south0_in00),
.o00(local0_out00),
.o01(east0_out00),
.o02(west0_out00),
.o03(north0_out00),
.o04(south0_out00)
);
router r001
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in01),
.i01(east0_in01),
.i02(west0_in01),
.i03(north0_in01),
.i04(south0_in01),
.o00(local0_out01),
.o01(east0_out01),
.o02(west0_out01),
.o03(north0_out01),
.o04(south0_out01)
);
router r002
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in02),
.i01(east0_in02),
.i02(west0_in02),
.i03(north0_in02),
.i04(south0_in02),
.o00(local0_out02),
.o01(east0_out02),
.o02(west0_out02),
.o03(north0_out02),
.o04(south0_out02)
);
router r003
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in03),
.i01(east0_in03),
.i02(west0_in03),
.i03(north0_in03),
.i04(south0_in03),
.o00(local0_out03),
.o01(east0_out03),
.o02(west0_out03),
.o03(north0_out03),
.o04(south0_out03)
);
router r004
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in04),
.i01(east0_in04),
.i02(west0_in04),
.i03(north0_in04),
.i04(south0_in04),
.o00(local0_out04),
.o01(east0_out04),
.o02(west0_out04),
.o03(north0_out04),
.o04(south0_out04)
);
router r005
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in05),
.i01(east0_in05),
.i02(west0_in05),
.i03(north0_in05),
.i04(south0_in05),
.o00(local0_out05),
.o01(east0_out05),
.o02(west0_out05),
.o03(north0_out05),
.o04(south0_out05)
);
router r006
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in06),
.i01(east0_in06),
.i02(west0_in06),
.i03(north0_in06),
.i04(south0_in06),
.o00(local0_out06),
.o01(east0_out06),
.o02(west0_out06),
.o03(north0_out06),
.o04(south0_out06)
);
router r007
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in07),
.i01(east0_in07),
.i02(west0_in07),
.i03(north0_in07),
.i04(south0_in07),
.o00(local0_out07),
.o01(east0_out07),
.o02(west0_out07),
.o03(north0_out07),
.o04(south0_out07)
);
router r008
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in08),
.i01(east0_in08),
.i02(west0_in08),
.i03(north0_in08),
.i04(south0_in08),
.o00(local0_out08),
.o01(east0_out08),
.o02(west0_out08),
.o03(north0_out08),
.o04(south0_out08)
);
router r009
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in09),
.i01(east0_in09),
.i02(west0_in09),
.i03(north0_in09),
.i04(south0_in09),
.o00(local0_out09),
.o01(east0_out09),
.o02(west0_out09),
.o03(north0_out09),
.o04(south0_out09)
);
router r0010
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in010),
.i01(east0_in010),
.i02(west0_in010),
.i03(north0_in010),
.i04(south0_in010),
.o00(local0_out010),
.o01(east0_out010),
.o02(west0_out010),
.o03(north0_out010),
.o04(south0_out010)
);
router r0011
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in011),
.i01(east0_in011),
.i02(west0_in011),
.i03(north0_in011),
.i04(south0_in011),
.o00(local0_out011),
.o01(east0_out011),
.o02(west0_out011),
.o03(north0_out011),
.o04(south0_out011)
);
router r0012
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in012),
.i01(east0_in012),
.i02(west0_in012),
.i03(north0_in012),
.i04(south0_in012),
.o00(local0_out012),
.o01(east0_out012),
.o02(west0_out012),
.o03(north0_out012),
.o04(south0_out012)
);
router r0013
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in013),
.i01(east0_in013),
.i02(west0_in013),
.i03(north0_in013),
.i04(south0_in013),
.o00(local0_out013),
.o01(east0_out013),
.o02(west0_out013),
.o03(north0_out013),
.o04(south0_out013)
);
router r0014
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in014),
.i01(east0_in014),
.i02(west0_in014),
.i03(north0_in014),
.i04(south0_in014),
.o00(local0_out014),
.o01(east0_out014),
.o02(west0_out014),
.o03(north0_out014),
.o04(south0_out014)
);
router r0015
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in015),
.i01(east0_in015),
.i02(west0_in015),
.i03(north0_in015),
.i04(south0_in015),
.o00(local0_out015),
.o01(east0_out015),
.o02(west0_out015),
.o03(north0_out015),
.o04(south0_out015)
);
router r110
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in10),
.i01(east1_in10),
.i02(west1_in10),
.i03(north1_in10),
.i04(south1_in10),
.o00(local1_out10),
.o01(east1_out10),
.o02(west1_out10),
.o03(north1_out10),
.o04(south1_out10)
);
router r111
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in11),
.i01(east1_in11),
.i02(west1_in11),
.i03(north1_in11),
.i04(south1_in11),
.o00(local1_out11),
.o01(east1_out11),
.o02(west1_out11),
.o03(north1_out11),
.o04(south1_out11)
);
router r112
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in12),
.i01(east1_in12),
.i02(west1_in12),
.i03(north1_in12),
.i04(south1_in12),
.o00(local1_out12),
.o01(east1_out12),
.o02(west1_out12),
.o03(north1_out12),
.o04(south1_out12)
);
router r113
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in13),
.i01(east1_in13),
.i02(west1_in13),
.i03(north1_in13),
.i04(south1_in13),
.o00(local1_out13),
.o01(east1_out13),
.o02(west1_out13),
.o03(north1_out13),
.o04(south1_out13)
);
router r114
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in14),
.i01(east1_in14),
.i02(west1_in14),
.i03(north1_in14),
.i04(south1_in14),
.o00(local1_out14),
.o01(east1_out14),
.o02(west1_out14),
.o03(north1_out14),
.o04(south1_out14)
);
router r115
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in15),
.i01(east1_in15),
.i02(west1_in15),
.i03(north1_in15),
.i04(south1_in15),
.o00(local1_out15),
.o01(east1_out15),
.o02(west1_out15),
.o03(north1_out15),
.o04(south1_out15)
);
router r116
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in16),
.i01(east1_in16),
.i02(west1_in16),
.i03(north1_in16),
.i04(south1_in16),
.o00(local1_out16),
.o01(east1_out16),
.o02(west1_out16),
.o03(north1_out16),
.o04(south1_out16)
);
router r117
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in17),
.i01(east1_in17),
.i02(west1_in17),
.i03(north1_in17),
.i04(south1_in17),
.o00(local1_out17),
.o01(east1_out17),
.o02(west1_out17),
.o03(north1_out17),
.o04(south1_out17)
);
router r118
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in18),
.i01(east1_in18),
.i02(west1_in18),
.i03(north1_in18),
.i04(south1_in18),
.o00(local1_out18),
.o01(east1_out18),
.o02(west1_out18),
.o03(north1_out18),
.o04(south1_out18)
);
router r119
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in19),
.i01(east1_in19),
.i02(west1_in19),
.i03(north1_in19),
.i04(south1_in19),
.o00(local1_out19),
.o01(east1_out19),
.o02(west1_out19),
.o03(north1_out19),
.o04(south1_out19)
);
router r1110
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in110),
.i01(east1_in110),
.i02(west1_in110),
.i03(north1_in110),
.i04(south1_in110),
.o00(local1_out110),
.o01(east1_out110),
.o02(west1_out110),
.o03(north1_out110),
.o04(south1_out110)
);
router r1111
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in111),
.i01(east1_in111),
.i02(west1_in111),
.i03(north1_in111),
.i04(south1_in111),
.o00(local1_out111),
.o01(east1_out111),
.o02(west1_out111),
.o03(north1_out111),
.o04(south1_out111)
);
router r1112
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in112),
.i01(east1_in112),
.i02(west1_in112),
.i03(north1_in112),
.i04(south1_in112),
.o00(local1_out112),
.o01(east1_out112),
.o02(west1_out112),
.o03(north1_out112),
.o04(south1_out112)
);
router r1113
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in113),
.i01(east1_in113),
.i02(west1_in113),
.i03(north1_in113),
.i04(south1_in113),
.o00(local1_out113),
.o01(east1_out113),
.o02(west1_out113),
.o03(north1_out113),
.o04(south1_out113)
);
router r1114
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in114),
.i01(east1_in114),
.i02(west1_in114),
.i03(north1_in114),
.i04(south1_in114),
.o00(local1_out114),
.o01(east1_out114),
.o02(west1_out114),
.o03(north1_out114),
.o04(south1_out114)
);
router r1115
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in115),
.i01(east1_in115),
.i02(west1_in115),
.i03(north1_in115),
.i04(south1_in115),
.o00(local1_out115),
.o01(east1_out115),
.o02(west1_out115),
.o03(north1_out115),
.o04(south1_out115)
);
router r220
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in20),
.i01(east2_in20),
.i02(west2_in20),
.i03(north2_in20),
.i04(south2_in20),
.o00(local2_out20),
.o01(east2_out20),
.o02(west2_out20),
.o03(north2_out20),
.o04(south2_out20)
);
router r221
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in21),
.i01(east2_in21),
.i02(west2_in21),
.i03(north2_in21),
.i04(south2_in21),
.o00(local2_out21),
.o01(east2_out21),
.o02(west2_out21),
.o03(north2_out21),
.o04(south2_out21)
);
router r222
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in22),
.i01(east2_in22),
.i02(west2_in22),
.i03(north2_in22),
.i04(south2_in22),
.o00(local2_out22),
.o01(east2_out22),
.o02(west2_out22),
.o03(north2_out22),
.o04(south2_out22)
);
router r223
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in23),
.i01(east2_in23),
.i02(west2_in23),
.i03(north2_in23),
.i04(south2_in23),
.o00(local2_out23),
.o01(east2_out23),
.o02(west2_out23),
.o03(north2_out23),
.o04(south2_out23)
);
router r224
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in24),
.i01(east2_in24),
.i02(west2_in24),
.i03(north2_in24),
.i04(south2_in24),
.o00(local2_out24),
.o01(east2_out24),
.o02(west2_out24),
.o03(north2_out24),
.o04(south2_out24)
);
router r225
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in25),
.i01(east2_in25),
.i02(west2_in25),
.i03(north2_in25),
.i04(south2_in25),
.o00(local2_out25),
.o01(east2_out25),
.o02(west2_out25),
.o03(north2_out25),
.o04(south2_out25)
);
router r226
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in26),
.i01(east2_in26),
.i02(west2_in26),
.i03(north2_in26),
.i04(south2_in26),
.o00(local2_out26),
.o01(east2_out26),
.o02(west2_out26),
.o03(north2_out26),
.o04(south2_out26)
);
router r227
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in27),
.i01(east2_in27),
.i02(west2_in27),
.i03(north2_in27),
.i04(south2_in27),
.o00(local2_out27),
.o01(east2_out27),
.o02(west2_out27),
.o03(north2_out27),
.o04(south2_out27)
);
router r228
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in28),
.i01(east2_in28),
.i02(west2_in28),
.i03(north2_in28),
.i04(south2_in28),
.o00(local2_out28),
.o01(east2_out28),
.o02(west2_out28),
.o03(north2_out28),
.o04(south2_out28)
);
router r229
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in29),
.i01(east2_in29),
.i02(west2_in29),
.i03(north2_in29),
.i04(south2_in29),
.o00(local2_out29),
.o01(east2_out29),
.o02(west2_out29),
.o03(north2_out29),
.o04(south2_out29)
);
router r2210
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in210),
.i01(east2_in210),
.i02(west2_in210),
.i03(north2_in210),
.i04(south2_in210),
.o00(local2_out210),
.o01(east2_out210),
.o02(west2_out210),
.o03(north2_out210),
.o04(south2_out210)
);
router r2211
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in211),
.i01(east2_in211),
.i02(west2_in211),
.i03(north2_in211),
.i04(south2_in211),
.o00(local2_out211),
.o01(east2_out211),
.o02(west2_out211),
.o03(north2_out211),
.o04(south2_out211)
);
router r2212
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in212),
.i01(east2_in212),
.i02(west2_in212),
.i03(north2_in212),
.i04(south2_in212),
.o00(local2_out212),
.o01(east2_out212),
.o02(west2_out212),
.o03(north2_out212),
.o04(south2_out212)
);
router r2213
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in213),
.i01(east2_in213),
.i02(west2_in213),
.i03(north2_in213),
.i04(south2_in213),
.o00(local2_out213),
.o01(east2_out213),
.o02(west2_out213),
.o03(north2_out213),
.o04(south2_out213)
);
router r2214
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in214),
.i01(east2_in214),
.i02(west2_in214),
.i03(north2_in214),
.i04(south2_in214),
.o00(local2_out214),
.o01(east2_out214),
.o02(west2_out214),
.o03(north2_out214),
.o04(south2_out214)
);
router r2215
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in215),
.i01(east2_in215),
.i02(west2_in215),
.i03(north2_in215),
.i04(south2_in215),
.o00(local2_out215),
.o01(east2_out215),
.o02(west2_out215),
.o03(north2_out215),
.o04(south2_out215)
);
router r330
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in30),
.i01(east3_in30),
.i02(west3_in30),
.i03(north3_in30),
.i04(south3_in30),
.o00(local3_out30),
.o01(east3_out30),
.o02(west3_out30),
.o03(north3_out30),
.o04(south3_out30)
);
router r331
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in31),
.i01(east3_in31),
.i02(west3_in31),
.i03(north3_in31),
.i04(south3_in31),
.o00(local3_out31),
.o01(east3_out31),
.o02(west3_out31),
.o03(north3_out31),
.o04(south3_out31)
);
router r332
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in32),
.i01(east3_in32),
.i02(west3_in32),
.i03(north3_in32),
.i04(south3_in32),
.o00(local3_out32),
.o01(east3_out32),
.o02(west3_out32),
.o03(north3_out32),
.o04(south3_out32)
);
router r333
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in33),
.i01(east3_in33),
.i02(west3_in33),
.i03(north3_in33),
.i04(south3_in33),
.o00(local3_out33),
.o01(east3_out33),
.o02(west3_out33),
.o03(north3_out33),
.o04(south3_out33)
);
router r334
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in34),
.i01(east3_in34),
.i02(west3_in34),
.i03(north3_in34),
.i04(south3_in34),
.o00(local3_out34),
.o01(east3_out34),
.o02(west3_out34),
.o03(north3_out34),
.o04(south3_out34)
);
router r335
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in35),
.i01(east3_in35),
.i02(west3_in35),
.i03(north3_in35),
.i04(south3_in35),
.o00(local3_out35),
.o01(east3_out35),
.o02(west3_out35),
.o03(north3_out35),
.o04(south3_out35)
);
router r336
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in36),
.i01(east3_in36),
.i02(west3_in36),
.i03(north3_in36),
.i04(south3_in36),
.o00(local3_out36),
.o01(east3_out36),
.o02(west3_out36),
.o03(north3_out36),
.o04(south3_out36)
);
router r337
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in37),
.i01(east3_in37),
.i02(west3_in37),
.i03(north3_in37),
.i04(south3_in37),
.o00(local3_out37),
.o01(east3_out37),
.o02(west3_out37),
.o03(north3_out37),
.o04(south3_out37)
);
router r338
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in38),
.i01(east3_in38),
.i02(west3_in38),
.i03(north3_in38),
.i04(south3_in38),
.o00(local3_out38),
.o01(east3_out38),
.o02(west3_out38),
.o03(north3_out38),
.o04(south3_out38)
);
router r339
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in39),
.i01(east3_in39),
.i02(west3_in39),
.i03(north3_in39),
.i04(south3_in39),
.o00(local3_out39),
.o01(east3_out39),
.o02(west3_out39),
.o03(north3_out39),
.o04(south3_out39)
);
router r3310
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in310),
.i01(east3_in310),
.i02(west3_in310),
.i03(north3_in310),
.i04(south3_in310),
.o00(local3_out310),
.o01(east3_out310),
.o02(west3_out310),
.o03(north3_out310),
.o04(south3_out310)
);
router r3311
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in311),
.i01(east3_in311),
.i02(west3_in311),
.i03(north3_in311),
.i04(south3_in311),
.o00(local3_out311),
.o01(east3_out311),
.o02(west3_out311),
.o03(north3_out311),
.o04(south3_out311)
);
router r3312
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in312),
.i01(east3_in312),
.i02(west3_in312),
.i03(north3_in312),
.i04(south3_in312),
.o00(local3_out312),
.o01(east3_out312),
.o02(west3_out312),
.o03(north3_out312),
.o04(south3_out312)
);
router r3313
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in313),
.i01(east3_in313),
.i02(west3_in313),
.i03(north3_in313),
.i04(south3_in313),
.o00(local3_out313),
.o01(east3_out313),
.o02(west3_out313),
.o03(north3_out313),
.o04(south3_out313)
);
router r3314
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in314),
.i01(east3_in314),
.i02(west3_in314),
.i03(north3_in314),
.i04(south3_in314),
.o00(local3_out314),
.o01(east3_out314),
.o02(west3_out314),
.o03(north3_out314),
.o04(south3_out314)
);
router r3315
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in315),
.i01(east3_in315),
.i02(west3_in315),
.i03(north3_in315),
.i04(south3_in315),
.o00(local3_out315),
.o01(east3_out315),
.o02(west3_out315),
.o03(north3_out315),
.o04(south3_out315)
);
router r440
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in40),
.i01(east4_in40),
.i02(west4_in40),
.i03(north4_in40),
.i04(south4_in40),
.o00(local4_out40),
.o01(east4_out40),
.o02(west4_out40),
.o03(north4_out40),
.o04(south4_out40)
);
router r441
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in41),
.i01(east4_in41),
.i02(west4_in41),
.i03(north4_in41),
.i04(south4_in41),
.o00(local4_out41),
.o01(east4_out41),
.o02(west4_out41),
.o03(north4_out41),
.o04(south4_out41)
);
router r442
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in42),
.i01(east4_in42),
.i02(west4_in42),
.i03(north4_in42),
.i04(south4_in42),
.o00(local4_out42),
.o01(east4_out42),
.o02(west4_out42),
.o03(north4_out42),
.o04(south4_out42)
);
router r443
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in43),
.i01(east4_in43),
.i02(west4_in43),
.i03(north4_in43),
.i04(south4_in43),
.o00(local4_out43),
.o01(east4_out43),
.o02(west4_out43),
.o03(north4_out43),
.o04(south4_out43)
);
router r444
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in44),
.i01(east4_in44),
.i02(west4_in44),
.i03(north4_in44),
.i04(south4_in44),
.o00(local4_out44),
.o01(east4_out44),
.o02(west4_out44),
.o03(north4_out44),
.o04(south4_out44)
);
router r445
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in45),
.i01(east4_in45),
.i02(west4_in45),
.i03(north4_in45),
.i04(south4_in45),
.o00(local4_out45),
.o01(east4_out45),
.o02(west4_out45),
.o03(north4_out45),
.o04(south4_out45)
);
router r446
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in46),
.i01(east4_in46),
.i02(west4_in46),
.i03(north4_in46),
.i04(south4_in46),
.o00(local4_out46),
.o01(east4_out46),
.o02(west4_out46),
.o03(north4_out46),
.o04(south4_out46)
);
router r447
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in47),
.i01(east4_in47),
.i02(west4_in47),
.i03(north4_in47),
.i04(south4_in47),
.o00(local4_out47),
.o01(east4_out47),
.o02(west4_out47),
.o03(north4_out47),
.o04(south4_out47)
);
router r448
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in48),
.i01(east4_in48),
.i02(west4_in48),
.i03(north4_in48),
.i04(south4_in48),
.o00(local4_out48),
.o01(east4_out48),
.o02(west4_out48),
.o03(north4_out48),
.o04(south4_out48)
);
router r449
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in49),
.i01(east4_in49),
.i02(west4_in49),
.i03(north4_in49),
.i04(south4_in49),
.o00(local4_out49),
.o01(east4_out49),
.o02(west4_out49),
.o03(north4_out49),
.o04(south4_out49)
);
router r4410
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in410),
.i01(east4_in410),
.i02(west4_in410),
.i03(north4_in410),
.i04(south4_in410),
.o00(local4_out410),
.o01(east4_out410),
.o02(west4_out410),
.o03(north4_out410),
.o04(south4_out410)
);
router r4411
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in411),
.i01(east4_in411),
.i02(west4_in411),
.i03(north4_in411),
.i04(south4_in411),
.o00(local4_out411),
.o01(east4_out411),
.o02(west4_out411),
.o03(north4_out411),
.o04(south4_out411)
);
router r4412
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in412),
.i01(east4_in412),
.i02(west4_in412),
.i03(north4_in412),
.i04(south4_in412),
.o00(local4_out412),
.o01(east4_out412),
.o02(west4_out412),
.o03(north4_out412),
.o04(south4_out412)
);
router r4413
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in413),
.i01(east4_in413),
.i02(west4_in413),
.i03(north4_in413),
.i04(south4_in413),
.o00(local4_out413),
.o01(east4_out413),
.o02(west4_out413),
.o03(north4_out413),
.o04(south4_out413)
);
router r4414
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in414),
.i01(east4_in414),
.i02(west4_in414),
.i03(north4_in414),
.i04(south4_in414),
.o00(local4_out414),
.o01(east4_out414),
.o02(west4_out414),
.o03(north4_out414),
.o04(south4_out414)
);
router r4415
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in415),
.i01(east4_in415),
.i02(west4_in415),
.i03(north4_in415),
.i04(south4_in415),
.o00(local4_out415),
.o01(east4_out415),
.o02(west4_out415),
.o03(north4_out415),
.o04(south4_out415)
);
router r550
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in50),
.i01(east5_in50),
.i02(west5_in50),
.i03(north5_in50),
.i04(south5_in50),
.o00(local5_out50),
.o01(east5_out50),
.o02(west5_out50),
.o03(north5_out50),
.o04(south5_out50)
);
router r551
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in51),
.i01(east5_in51),
.i02(west5_in51),
.i03(north5_in51),
.i04(south5_in51),
.o00(local5_out51),
.o01(east5_out51),
.o02(west5_out51),
.o03(north5_out51),
.o04(south5_out51)
);
router r552
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in52),
.i01(east5_in52),
.i02(west5_in52),
.i03(north5_in52),
.i04(south5_in52),
.o00(local5_out52),
.o01(east5_out52),
.o02(west5_out52),
.o03(north5_out52),
.o04(south5_out52)
);
router r553
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in53),
.i01(east5_in53),
.i02(west5_in53),
.i03(north5_in53),
.i04(south5_in53),
.o00(local5_out53),
.o01(east5_out53),
.o02(west5_out53),
.o03(north5_out53),
.o04(south5_out53)
);
router r554
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in54),
.i01(east5_in54),
.i02(west5_in54),
.i03(north5_in54),
.i04(south5_in54),
.o00(local5_out54),
.o01(east5_out54),
.o02(west5_out54),
.o03(north5_out54),
.o04(south5_out54)
);
router r555
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in55),
.i01(east5_in55),
.i02(west5_in55),
.i03(north5_in55),
.i04(south5_in55),
.o00(local5_out55),
.o01(east5_out55),
.o02(west5_out55),
.o03(north5_out55),
.o04(south5_out55)
);
router r556
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in56),
.i01(east5_in56),
.i02(west5_in56),
.i03(north5_in56),
.i04(south5_in56),
.o00(local5_out56),
.o01(east5_out56),
.o02(west5_out56),
.o03(north5_out56),
.o04(south5_out56)
);
router r557
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in57),
.i01(east5_in57),
.i02(west5_in57),
.i03(north5_in57),
.i04(south5_in57),
.o00(local5_out57),
.o01(east5_out57),
.o02(west5_out57),
.o03(north5_out57),
.o04(south5_out57)
);
router r558
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in58),
.i01(east5_in58),
.i02(west5_in58),
.i03(north5_in58),
.i04(south5_in58),
.o00(local5_out58),
.o01(east5_out58),
.o02(west5_out58),
.o03(north5_out58),
.o04(south5_out58)
);
router r559
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in59),
.i01(east5_in59),
.i02(west5_in59),
.i03(north5_in59),
.i04(south5_in59),
.o00(local5_out59),
.o01(east5_out59),
.o02(west5_out59),
.o03(north5_out59),
.o04(south5_out59)
);
router r5510
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in510),
.i01(east5_in510),
.i02(west5_in510),
.i03(north5_in510),
.i04(south5_in510),
.o00(local5_out510),
.o01(east5_out510),
.o02(west5_out510),
.o03(north5_out510),
.o04(south5_out510)
);
router r5511
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in511),
.i01(east5_in511),
.i02(west5_in511),
.i03(north5_in511),
.i04(south5_in511),
.o00(local5_out511),
.o01(east5_out511),
.o02(west5_out511),
.o03(north5_out511),
.o04(south5_out511)
);
router r5512
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in512),
.i01(east5_in512),
.i02(west5_in512),
.i03(north5_in512),
.i04(south5_in512),
.o00(local5_out512),
.o01(east5_out512),
.o02(west5_out512),
.o03(north5_out512),
.o04(south5_out512)
);
router r5513
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in513),
.i01(east5_in513),
.i02(west5_in513),
.i03(north5_in513),
.i04(south5_in513),
.o00(local5_out513),
.o01(east5_out513),
.o02(west5_out513),
.o03(north5_out513),
.o04(south5_out513)
);
router r5514
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in514),
.i01(east5_in514),
.i02(west5_in514),
.i03(north5_in514),
.i04(south5_in514),
.o00(local5_out514),
.o01(east5_out514),
.o02(west5_out514),
.o03(north5_out514),
.o04(south5_out514)
);
router r5515
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in515),
.i01(east5_in515),
.i02(west5_in515),
.i03(north5_in515),
.i04(south5_in515),
.o00(local5_out515),
.o01(east5_out515),
.o02(west5_out515),
.o03(north5_out515),
.o04(south5_out515)
);
router r660
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in60),
.i01(east6_in60),
.i02(west6_in60),
.i03(north6_in60),
.i04(south6_in60),
.o00(local6_out60),
.o01(east6_out60),
.o02(west6_out60),
.o03(north6_out60),
.o04(south6_out60)
);
router r661
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in61),
.i01(east6_in61),
.i02(west6_in61),
.i03(north6_in61),
.i04(south6_in61),
.o00(local6_out61),
.o01(east6_out61),
.o02(west6_out61),
.o03(north6_out61),
.o04(south6_out61)
);
router r662
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in62),
.i01(east6_in62),
.i02(west6_in62),
.i03(north6_in62),
.i04(south6_in62),
.o00(local6_out62),
.o01(east6_out62),
.o02(west6_out62),
.o03(north6_out62),
.o04(south6_out62)
);
router r663
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in63),
.i01(east6_in63),
.i02(west6_in63),
.i03(north6_in63),
.i04(south6_in63),
.o00(local6_out63),
.o01(east6_out63),
.o02(west6_out63),
.o03(north6_out63),
.o04(south6_out63)
);
router r664
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in64),
.i01(east6_in64),
.i02(west6_in64),
.i03(north6_in64),
.i04(south6_in64),
.o00(local6_out64),
.o01(east6_out64),
.o02(west6_out64),
.o03(north6_out64),
.o04(south6_out64)
);
router r665
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in65),
.i01(east6_in65),
.i02(west6_in65),
.i03(north6_in65),
.i04(south6_in65),
.o00(local6_out65),
.o01(east6_out65),
.o02(west6_out65),
.o03(north6_out65),
.o04(south6_out65)
);
router r666
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in66),
.i01(east6_in66),
.i02(west6_in66),
.i03(north6_in66),
.i04(south6_in66),
.o00(local6_out66),
.o01(east6_out66),
.o02(west6_out66),
.o03(north6_out66),
.o04(south6_out66)
);
router r667
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in67),
.i01(east6_in67),
.i02(west6_in67),
.i03(north6_in67),
.i04(south6_in67),
.o00(local6_out67),
.o01(east6_out67),
.o02(west6_out67),
.o03(north6_out67),
.o04(south6_out67)
);
router r668
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in68),
.i01(east6_in68),
.i02(west6_in68),
.i03(north6_in68),
.i04(south6_in68),
.o00(local6_out68),
.o01(east6_out68),
.o02(west6_out68),
.o03(north6_out68),
.o04(south6_out68)
);
router r669
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in69),
.i01(east6_in69),
.i02(west6_in69),
.i03(north6_in69),
.i04(south6_in69),
.o00(local6_out69),
.o01(east6_out69),
.o02(west6_out69),
.o03(north6_out69),
.o04(south6_out69)
);
router r6610
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in610),
.i01(east6_in610),
.i02(west6_in610),
.i03(north6_in610),
.i04(south6_in610),
.o00(local6_out610),
.o01(east6_out610),
.o02(west6_out610),
.o03(north6_out610),
.o04(south6_out610)
);
router r6611
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in611),
.i01(east6_in611),
.i02(west6_in611),
.i03(north6_in611),
.i04(south6_in611),
.o00(local6_out611),
.o01(east6_out611),
.o02(west6_out611),
.o03(north6_out611),
.o04(south6_out611)
);
router r6612
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in612),
.i01(east6_in612),
.i02(west6_in612),
.i03(north6_in612),
.i04(south6_in612),
.o00(local6_out612),
.o01(east6_out612),
.o02(west6_out612),
.o03(north6_out612),
.o04(south6_out612)
);
router r6613
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in613),
.i01(east6_in613),
.i02(west6_in613),
.i03(north6_in613),
.i04(south6_in613),
.o00(local6_out613),
.o01(east6_out613),
.o02(west6_out613),
.o03(north6_out613),
.o04(south6_out613)
);
router r6614
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in614),
.i01(east6_in614),
.i02(west6_in614),
.i03(north6_in614),
.i04(south6_in614),
.o00(local6_out614),
.o01(east6_out614),
.o02(west6_out614),
.o03(north6_out614),
.o04(south6_out614)
);
router r6615
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in615),
.i01(east6_in615),
.i02(west6_in615),
.i03(north6_in615),
.i04(south6_in615),
.o00(local6_out615),
.o01(east6_out615),
.o02(west6_out615),
.o03(north6_out615),
.o04(south6_out615)
);
router r770
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in70),
.i01(east7_in70),
.i02(west7_in70),
.i03(north7_in70),
.i04(south7_in70),
.o00(local7_out70),
.o01(east7_out70),
.o02(west7_out70),
.o03(north7_out70),
.o04(south7_out70)
);
router r771
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in71),
.i01(east7_in71),
.i02(west7_in71),
.i03(north7_in71),
.i04(south7_in71),
.o00(local7_out71),
.o01(east7_out71),
.o02(west7_out71),
.o03(north7_out71),
.o04(south7_out71)
);
router r772
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in72),
.i01(east7_in72),
.i02(west7_in72),
.i03(north7_in72),
.i04(south7_in72),
.o00(local7_out72),
.o01(east7_out72),
.o02(west7_out72),
.o03(north7_out72),
.o04(south7_out72)
);
router r773
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in73),
.i01(east7_in73),
.i02(west7_in73),
.i03(north7_in73),
.i04(south7_in73),
.o00(local7_out73),
.o01(east7_out73),
.o02(west7_out73),
.o03(north7_out73),
.o04(south7_out73)
);
router r774
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in74),
.i01(east7_in74),
.i02(west7_in74),
.i03(north7_in74),
.i04(south7_in74),
.o00(local7_out74),
.o01(east7_out74),
.o02(west7_out74),
.o03(north7_out74),
.o04(south7_out74)
);
router r775
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in75),
.i01(east7_in75),
.i02(west7_in75),
.i03(north7_in75),
.i04(south7_in75),
.o00(local7_out75),
.o01(east7_out75),
.o02(west7_out75),
.o03(north7_out75),
.o04(south7_out75)
);
router r776
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in76),
.i01(east7_in76),
.i02(west7_in76),
.i03(north7_in76),
.i04(south7_in76),
.o00(local7_out76),
.o01(east7_out76),
.o02(west7_out76),
.o03(north7_out76),
.o04(south7_out76)
);
router r777
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in77),
.i01(east7_in77),
.i02(west7_in77),
.i03(north7_in77),
.i04(south7_in77),
.o00(local7_out77),
.o01(east7_out77),
.o02(west7_out77),
.o03(north7_out77),
.o04(south7_out77)
);
router r778
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in78),
.i01(east7_in78),
.i02(west7_in78),
.i03(north7_in78),
.i04(south7_in78),
.o00(local7_out78),
.o01(east7_out78),
.o02(west7_out78),
.o03(north7_out78),
.o04(south7_out78)
);
router r779
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in79),
.i01(east7_in79),
.i02(west7_in79),
.i03(north7_in79),
.i04(south7_in79),
.o00(local7_out79),
.o01(east7_out79),
.o02(west7_out79),
.o03(north7_out79),
.o04(south7_out79)
);
router r7710
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in710),
.i01(east7_in710),
.i02(west7_in710),
.i03(north7_in710),
.i04(south7_in710),
.o00(local7_out710),
.o01(east7_out710),
.o02(west7_out710),
.o03(north7_out710),
.o04(south7_out710)
);
router r7711
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in711),
.i01(east7_in711),
.i02(west7_in711),
.i03(north7_in711),
.i04(south7_in711),
.o00(local7_out711),
.o01(east7_out711),
.o02(west7_out711),
.o03(north7_out711),
.o04(south7_out711)
);
router r7712
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in712),
.i01(east7_in712),
.i02(west7_in712),
.i03(north7_in712),
.i04(south7_in712),
.o00(local7_out712),
.o01(east7_out712),
.o02(west7_out712),
.o03(north7_out712),
.o04(south7_out712)
);
router r7713
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in713),
.i01(east7_in713),
.i02(west7_in713),
.i03(north7_in713),
.i04(south7_in713),
.o00(local7_out713),
.o01(east7_out713),
.o02(west7_out713),
.o03(north7_out713),
.o04(south7_out713)
);
router r7714
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in714),
.i01(east7_in714),
.i02(west7_in714),
.i03(north7_in714),
.i04(south7_in714),
.o00(local7_out714),
.o01(east7_out714),
.o02(west7_out714),
.o03(north7_out714),
.o04(south7_out714)
);
router r7715
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in715),
.i01(east7_in715),
.i02(west7_in715),
.i03(north7_in715),
.i04(south7_in715),
.o00(local7_out715),
.o01(east7_out715),
.o02(west7_out715),
.o03(north7_out715),
.o04(south7_out715)
);
router r880
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in80),
.i01(east8_in80),
.i02(west8_in80),
.i03(north8_in80),
.i04(south8_in80),
.o00(local8_out80),
.o01(east8_out80),
.o02(west8_out80),
.o03(north8_out80),
.o04(south8_out80)
);
router r881
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in81),
.i01(east8_in81),
.i02(west8_in81),
.i03(north8_in81),
.i04(south8_in81),
.o00(local8_out81),
.o01(east8_out81),
.o02(west8_out81),
.o03(north8_out81),
.o04(south8_out81)
);
router r882
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in82),
.i01(east8_in82),
.i02(west8_in82),
.i03(north8_in82),
.i04(south8_in82),
.o00(local8_out82),
.o01(east8_out82),
.o02(west8_out82),
.o03(north8_out82),
.o04(south8_out82)
);
router r883
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in83),
.i01(east8_in83),
.i02(west8_in83),
.i03(north8_in83),
.i04(south8_in83),
.o00(local8_out83),
.o01(east8_out83),
.o02(west8_out83),
.o03(north8_out83),
.o04(south8_out83)
);
router r884
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in84),
.i01(east8_in84),
.i02(west8_in84),
.i03(north8_in84),
.i04(south8_in84),
.o00(local8_out84),
.o01(east8_out84),
.o02(west8_out84),
.o03(north8_out84),
.o04(south8_out84)
);
router r885
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in85),
.i01(east8_in85),
.i02(west8_in85),
.i03(north8_in85),
.i04(south8_in85),
.o00(local8_out85),
.o01(east8_out85),
.o02(west8_out85),
.o03(north8_out85),
.o04(south8_out85)
);
router r886
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in86),
.i01(east8_in86),
.i02(west8_in86),
.i03(north8_in86),
.i04(south8_in86),
.o00(local8_out86),
.o01(east8_out86),
.o02(west8_out86),
.o03(north8_out86),
.o04(south8_out86)
);
router r887
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in87),
.i01(east8_in87),
.i02(west8_in87),
.i03(north8_in87),
.i04(south8_in87),
.o00(local8_out87),
.o01(east8_out87),
.o02(west8_out87),
.o03(north8_out87),
.o04(south8_out87)
);
router r888
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in88),
.i01(east8_in88),
.i02(west8_in88),
.i03(north8_in88),
.i04(south8_in88),
.o00(local8_out88),
.o01(east8_out88),
.o02(west8_out88),
.o03(north8_out88),
.o04(south8_out88)
);
router r889
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in89),
.i01(east8_in89),
.i02(west8_in89),
.i03(north8_in89),
.i04(south8_in89),
.o00(local8_out89),
.o01(east8_out89),
.o02(west8_out89),
.o03(north8_out89),
.o04(south8_out89)
);
router r8810
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in810),
.i01(east8_in810),
.i02(west8_in810),
.i03(north8_in810),
.i04(south8_in810),
.o00(local8_out810),
.o01(east8_out810),
.o02(west8_out810),
.o03(north8_out810),
.o04(south8_out810)
);
router r8811
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in811),
.i01(east8_in811),
.i02(west8_in811),
.i03(north8_in811),
.i04(south8_in811),
.o00(local8_out811),
.o01(east8_out811),
.o02(west8_out811),
.o03(north8_out811),
.o04(south8_out811)
);
router r8812
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in812),
.i01(east8_in812),
.i02(west8_in812),
.i03(north8_in812),
.i04(south8_in812),
.o00(local8_out812),
.o01(east8_out812),
.o02(west8_out812),
.o03(north8_out812),
.o04(south8_out812)
);
router r8813
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in813),
.i01(east8_in813),
.i02(west8_in813),
.i03(north8_in813),
.i04(south8_in813),
.o00(local8_out813),
.o01(east8_out813),
.o02(west8_out813),
.o03(north8_out813),
.o04(south8_out813)
);
router r8814
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in814),
.i01(east8_in814),
.i02(west8_in814),
.i03(north8_in814),
.i04(south8_in814),
.o00(local8_out814),
.o01(east8_out814),
.o02(west8_out814),
.o03(north8_out814),
.o04(south8_out814)
);
router r8815
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in815),
.i01(east8_in815),
.i02(west8_in815),
.i03(north8_in815),
.i04(south8_in815),
.o00(local8_out815),
.o01(east8_out815),
.o02(west8_out815),
.o03(north8_out815),
.o04(south8_out815)
);
router r990
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in90),
.i01(east9_in90),
.i02(west9_in90),
.i03(north9_in90),
.i04(south9_in90),
.o00(local9_out90),
.o01(east9_out90),
.o02(west9_out90),
.o03(north9_out90),
.o04(south9_out90)
);
router r991
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in91),
.i01(east9_in91),
.i02(west9_in91),
.i03(north9_in91),
.i04(south9_in91),
.o00(local9_out91),
.o01(east9_out91),
.o02(west9_out91),
.o03(north9_out91),
.o04(south9_out91)
);
router r992
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in92),
.i01(east9_in92),
.i02(west9_in92),
.i03(north9_in92),
.i04(south9_in92),
.o00(local9_out92),
.o01(east9_out92),
.o02(west9_out92),
.o03(north9_out92),
.o04(south9_out92)
);
router r993
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in93),
.i01(east9_in93),
.i02(west9_in93),
.i03(north9_in93),
.i04(south9_in93),
.o00(local9_out93),
.o01(east9_out93),
.o02(west9_out93),
.o03(north9_out93),
.o04(south9_out93)
);
router r994
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in94),
.i01(east9_in94),
.i02(west9_in94),
.i03(north9_in94),
.i04(south9_in94),
.o00(local9_out94),
.o01(east9_out94),
.o02(west9_out94),
.o03(north9_out94),
.o04(south9_out94)
);
router r995
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in95),
.i01(east9_in95),
.i02(west9_in95),
.i03(north9_in95),
.i04(south9_in95),
.o00(local9_out95),
.o01(east9_out95),
.o02(west9_out95),
.o03(north9_out95),
.o04(south9_out95)
);
router r996
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in96),
.i01(east9_in96),
.i02(west9_in96),
.i03(north9_in96),
.i04(south9_in96),
.o00(local9_out96),
.o01(east9_out96),
.o02(west9_out96),
.o03(north9_out96),
.o04(south9_out96)
);
router r997
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in97),
.i01(east9_in97),
.i02(west9_in97),
.i03(north9_in97),
.i04(south9_in97),
.o00(local9_out97),
.o01(east9_out97),
.o02(west9_out97),
.o03(north9_out97),
.o04(south9_out97)
);
router r998
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in98),
.i01(east9_in98),
.i02(west9_in98),
.i03(north9_in98),
.i04(south9_in98),
.o00(local9_out98),
.o01(east9_out98),
.o02(west9_out98),
.o03(north9_out98),
.o04(south9_out98)
);
router r999
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in99),
.i01(east9_in99),
.i02(west9_in99),
.i03(north9_in99),
.i04(south9_in99),
.o00(local9_out99),
.o01(east9_out99),
.o02(west9_out99),
.o03(north9_out99),
.o04(south9_out99)
);
router r9910
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in910),
.i01(east9_in910),
.i02(west9_in910),
.i03(north9_in910),
.i04(south9_in910),
.o00(local9_out910),
.o01(east9_out910),
.o02(west9_out910),
.o03(north9_out910),
.o04(south9_out910)
);
router r9911
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in911),
.i01(east9_in911),
.i02(west9_in911),
.i03(north9_in911),
.i04(south9_in911),
.o00(local9_out911),
.o01(east9_out911),
.o02(west9_out911),
.o03(north9_out911),
.o04(south9_out911)
);
router r9912
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in912),
.i01(east9_in912),
.i02(west9_in912),
.i03(north9_in912),
.i04(south9_in912),
.o00(local9_out912),
.o01(east9_out912),
.o02(west9_out912),
.o03(north9_out912),
.o04(south9_out912)
);
router r9913
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in913),
.i01(east9_in913),
.i02(west9_in913),
.i03(north9_in913),
.i04(south9_in913),
.o00(local9_out913),
.o01(east9_out913),
.o02(west9_out913),
.o03(north9_out913),
.o04(south9_out913)
);
router r9914
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in914),
.i01(east9_in914),
.i02(west9_in914),
.i03(north9_in914),
.i04(south9_in914),
.o00(local9_out914),
.o01(east9_out914),
.o02(west9_out914),
.o03(north9_out914),
.o04(south9_out914)
);
router r9915
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in915),
.i01(east9_in915),
.i02(west9_in915),
.i03(north9_in915),
.i04(south9_in915),
.o00(local9_out915),
.o01(east9_out915),
.o02(west9_out915),
.o03(north9_out915),
.o04(south9_out915)
);
router r10100
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in100),
.i01(east10_in100),
.i02(west10_in100),
.i03(north10_in100),
.i04(south10_in100),
.o00(local10_out100),
.o01(east10_out100),
.o02(west10_out100),
.o03(north10_out100),
.o04(south10_out100)
);
router r10101
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in101),
.i01(east10_in101),
.i02(west10_in101),
.i03(north10_in101),
.i04(south10_in101),
.o00(local10_out101),
.o01(east10_out101),
.o02(west10_out101),
.o03(north10_out101),
.o04(south10_out101)
);
router r10102
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in102),
.i01(east10_in102),
.i02(west10_in102),
.i03(north10_in102),
.i04(south10_in102),
.o00(local10_out102),
.o01(east10_out102),
.o02(west10_out102),
.o03(north10_out102),
.o04(south10_out102)
);
router r10103
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in103),
.i01(east10_in103),
.i02(west10_in103),
.i03(north10_in103),
.i04(south10_in103),
.o00(local10_out103),
.o01(east10_out103),
.o02(west10_out103),
.o03(north10_out103),
.o04(south10_out103)
);
router r10104
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in104),
.i01(east10_in104),
.i02(west10_in104),
.i03(north10_in104),
.i04(south10_in104),
.o00(local10_out104),
.o01(east10_out104),
.o02(west10_out104),
.o03(north10_out104),
.o04(south10_out104)
);
router r10105
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in105),
.i01(east10_in105),
.i02(west10_in105),
.i03(north10_in105),
.i04(south10_in105),
.o00(local10_out105),
.o01(east10_out105),
.o02(west10_out105),
.o03(north10_out105),
.o04(south10_out105)
);
router r10106
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in106),
.i01(east10_in106),
.i02(west10_in106),
.i03(north10_in106),
.i04(south10_in106),
.o00(local10_out106),
.o01(east10_out106),
.o02(west10_out106),
.o03(north10_out106),
.o04(south10_out106)
);
router r10107
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in107),
.i01(east10_in107),
.i02(west10_in107),
.i03(north10_in107),
.i04(south10_in107),
.o00(local10_out107),
.o01(east10_out107),
.o02(west10_out107),
.o03(north10_out107),
.o04(south10_out107)
);
router r10108
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in108),
.i01(east10_in108),
.i02(west10_in108),
.i03(north10_in108),
.i04(south10_in108),
.o00(local10_out108),
.o01(east10_out108),
.o02(west10_out108),
.o03(north10_out108),
.o04(south10_out108)
);
router r10109
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in109),
.i01(east10_in109),
.i02(west10_in109),
.i03(north10_in109),
.i04(south10_in109),
.o00(local10_out109),
.o01(east10_out109),
.o02(west10_out109),
.o03(north10_out109),
.o04(south10_out109)
);
router r101010
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in1010),
.i01(east10_in1010),
.i02(west10_in1010),
.i03(north10_in1010),
.i04(south10_in1010),
.o00(local10_out1010),
.o01(east10_out1010),
.o02(west10_out1010),
.o03(north10_out1010),
.o04(south10_out1010)
);
router r101011
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in1011),
.i01(east10_in1011),
.i02(west10_in1011),
.i03(north10_in1011),
.i04(south10_in1011),
.o00(local10_out1011),
.o01(east10_out1011),
.o02(west10_out1011),
.o03(north10_out1011),
.o04(south10_out1011)
);
router r101012
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in1012),
.i01(east10_in1012),
.i02(west10_in1012),
.i03(north10_in1012),
.i04(south10_in1012),
.o00(local10_out1012),
.o01(east10_out1012),
.o02(west10_out1012),
.o03(north10_out1012),
.o04(south10_out1012)
);
router r101013
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in1013),
.i01(east10_in1013),
.i02(west10_in1013),
.i03(north10_in1013),
.i04(south10_in1013),
.o00(local10_out1013),
.o01(east10_out1013),
.o02(west10_out1013),
.o03(north10_out1013),
.o04(south10_out1013)
);
router r101014
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in1014),
.i01(east10_in1014),
.i02(west10_in1014),
.i03(north10_in1014),
.i04(south10_in1014),
.o00(local10_out1014),
.o01(east10_out1014),
.o02(west10_out1014),
.o03(north10_out1014),
.o04(south10_out1014)
);
router r101015
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in1015),
.i01(east10_in1015),
.i02(west10_in1015),
.i03(north10_in1015),
.i04(south10_in1015),
.o00(local10_out1015),
.o01(east10_out1015),
.o02(west10_out1015),
.o03(north10_out1015),
.o04(south10_out1015)
);
router r11110
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in110),
.i01(east11_in110),
.i02(west11_in110),
.i03(north11_in110),
.i04(south11_in110),
.o00(local11_out110),
.o01(east11_out110),
.o02(west11_out110),
.o03(north11_out110),
.o04(south11_out110)
);
router r11111
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in111),
.i01(east11_in111),
.i02(west11_in111),
.i03(north11_in111),
.i04(south11_in111),
.o00(local11_out111),
.o01(east11_out111),
.o02(west11_out111),
.o03(north11_out111),
.o04(south11_out111)
);
router r11112
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in112),
.i01(east11_in112),
.i02(west11_in112),
.i03(north11_in112),
.i04(south11_in112),
.o00(local11_out112),
.o01(east11_out112),
.o02(west11_out112),
.o03(north11_out112),
.o04(south11_out112)
);
router r11113
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in113),
.i01(east11_in113),
.i02(west11_in113),
.i03(north11_in113),
.i04(south11_in113),
.o00(local11_out113),
.o01(east11_out113),
.o02(west11_out113),
.o03(north11_out113),
.o04(south11_out113)
);
router r11114
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in114),
.i01(east11_in114),
.i02(west11_in114),
.i03(north11_in114),
.i04(south11_in114),
.o00(local11_out114),
.o01(east11_out114),
.o02(west11_out114),
.o03(north11_out114),
.o04(south11_out114)
);
router r11115
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in115),
.i01(east11_in115),
.i02(west11_in115),
.i03(north11_in115),
.i04(south11_in115),
.o00(local11_out115),
.o01(east11_out115),
.o02(west11_out115),
.o03(north11_out115),
.o04(south11_out115)
);
router r11116
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in116),
.i01(east11_in116),
.i02(west11_in116),
.i03(north11_in116),
.i04(south11_in116),
.o00(local11_out116),
.o01(east11_out116),
.o02(west11_out116),
.o03(north11_out116),
.o04(south11_out116)
);
router r11117
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in117),
.i01(east11_in117),
.i02(west11_in117),
.i03(north11_in117),
.i04(south11_in117),
.o00(local11_out117),
.o01(east11_out117),
.o02(west11_out117),
.o03(north11_out117),
.o04(south11_out117)
);
router r11118
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in118),
.i01(east11_in118),
.i02(west11_in118),
.i03(north11_in118),
.i04(south11_in118),
.o00(local11_out118),
.o01(east11_out118),
.o02(west11_out118),
.o03(north11_out118),
.o04(south11_out118)
);
router r11119
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in119),
.i01(east11_in119),
.i02(west11_in119),
.i03(north11_in119),
.i04(south11_in119),
.o00(local11_out119),
.o01(east11_out119),
.o02(west11_out119),
.o03(north11_out119),
.o04(south11_out119)
);
router r111110
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in1110),
.i01(east11_in1110),
.i02(west11_in1110),
.i03(north11_in1110),
.i04(south11_in1110),
.o00(local11_out1110),
.o01(east11_out1110),
.o02(west11_out1110),
.o03(north11_out1110),
.o04(south11_out1110)
);
router r111111
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in1111),
.i01(east11_in1111),
.i02(west11_in1111),
.i03(north11_in1111),
.i04(south11_in1111),
.o00(local11_out1111),
.o01(east11_out1111),
.o02(west11_out1111),
.o03(north11_out1111),
.o04(south11_out1111)
);
router r111112
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in1112),
.i01(east11_in1112),
.i02(west11_in1112),
.i03(north11_in1112),
.i04(south11_in1112),
.o00(local11_out1112),
.o01(east11_out1112),
.o02(west11_out1112),
.o03(north11_out1112),
.o04(south11_out1112)
);
router r111113
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in1113),
.i01(east11_in1113),
.i02(west11_in1113),
.i03(north11_in1113),
.i04(south11_in1113),
.o00(local11_out1113),
.o01(east11_out1113),
.o02(west11_out1113),
.o03(north11_out1113),
.o04(south11_out1113)
);
router r111114
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in1114),
.i01(east11_in1114),
.i02(west11_in1114),
.i03(north11_in1114),
.i04(south11_in1114),
.o00(local11_out1114),
.o01(east11_out1114),
.o02(west11_out1114),
.o03(north11_out1114),
.o04(south11_out1114)
);
router r111115
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in1115),
.i01(east11_in1115),
.i02(west11_in1115),
.i03(north11_in1115),
.i04(south11_in1115),
.o00(local11_out1115),
.o01(east11_out1115),
.o02(west11_out1115),
.o03(north11_out1115),
.o04(south11_out1115)
);
router r12120
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in120),
.i01(east12_in120),
.i02(west12_in120),
.i03(north12_in120),
.i04(south12_in120),
.o00(local12_out120),
.o01(east12_out120),
.o02(west12_out120),
.o03(north12_out120),
.o04(south12_out120)
);
router r12121
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in121),
.i01(east12_in121),
.i02(west12_in121),
.i03(north12_in121),
.i04(south12_in121),
.o00(local12_out121),
.o01(east12_out121),
.o02(west12_out121),
.o03(north12_out121),
.o04(south12_out121)
);
router r12122
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in122),
.i01(east12_in122),
.i02(west12_in122),
.i03(north12_in122),
.i04(south12_in122),
.o00(local12_out122),
.o01(east12_out122),
.o02(west12_out122),
.o03(north12_out122),
.o04(south12_out122)
);
router r12123
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in123),
.i01(east12_in123),
.i02(west12_in123),
.i03(north12_in123),
.i04(south12_in123),
.o00(local12_out123),
.o01(east12_out123),
.o02(west12_out123),
.o03(north12_out123),
.o04(south12_out123)
);
router r12124
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in124),
.i01(east12_in124),
.i02(west12_in124),
.i03(north12_in124),
.i04(south12_in124),
.o00(local12_out124),
.o01(east12_out124),
.o02(west12_out124),
.o03(north12_out124),
.o04(south12_out124)
);
router r12125
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in125),
.i01(east12_in125),
.i02(west12_in125),
.i03(north12_in125),
.i04(south12_in125),
.o00(local12_out125),
.o01(east12_out125),
.o02(west12_out125),
.o03(north12_out125),
.o04(south12_out125)
);
router r12126
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in126),
.i01(east12_in126),
.i02(west12_in126),
.i03(north12_in126),
.i04(south12_in126),
.o00(local12_out126),
.o01(east12_out126),
.o02(west12_out126),
.o03(north12_out126),
.o04(south12_out126)
);
router r12127
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in127),
.i01(east12_in127),
.i02(west12_in127),
.i03(north12_in127),
.i04(south12_in127),
.o00(local12_out127),
.o01(east12_out127),
.o02(west12_out127),
.o03(north12_out127),
.o04(south12_out127)
);
router r12128
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in128),
.i01(east12_in128),
.i02(west12_in128),
.i03(north12_in128),
.i04(south12_in128),
.o00(local12_out128),
.o01(east12_out128),
.o02(west12_out128),
.o03(north12_out128),
.o04(south12_out128)
);
router r12129
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in129),
.i01(east12_in129),
.i02(west12_in129),
.i03(north12_in129),
.i04(south12_in129),
.o00(local12_out129),
.o01(east12_out129),
.o02(west12_out129),
.o03(north12_out129),
.o04(south12_out129)
);
router r121210
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in1210),
.i01(east12_in1210),
.i02(west12_in1210),
.i03(north12_in1210),
.i04(south12_in1210),
.o00(local12_out1210),
.o01(east12_out1210),
.o02(west12_out1210),
.o03(north12_out1210),
.o04(south12_out1210)
);
router r121211
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in1211),
.i01(east12_in1211),
.i02(west12_in1211),
.i03(north12_in1211),
.i04(south12_in1211),
.o00(local12_out1211),
.o01(east12_out1211),
.o02(west12_out1211),
.o03(north12_out1211),
.o04(south12_out1211)
);
router r121212
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in1212),
.i01(east12_in1212),
.i02(west12_in1212),
.i03(north12_in1212),
.i04(south12_in1212),
.o00(local12_out1212),
.o01(east12_out1212),
.o02(west12_out1212),
.o03(north12_out1212),
.o04(south12_out1212)
);
router r121213
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in1213),
.i01(east12_in1213),
.i02(west12_in1213),
.i03(north12_in1213),
.i04(south12_in1213),
.o00(local12_out1213),
.o01(east12_out1213),
.o02(west12_out1213),
.o03(north12_out1213),
.o04(south12_out1213)
);
router r121214
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in1214),
.i01(east12_in1214),
.i02(west12_in1214),
.i03(north12_in1214),
.i04(south12_in1214),
.o00(local12_out1214),
.o01(east12_out1214),
.o02(west12_out1214),
.o03(north12_out1214),
.o04(south12_out1214)
);
router r121215
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in1215),
.i01(east12_in1215),
.i02(west12_in1215),
.i03(north12_in1215),
.i04(south12_in1215),
.o00(local12_out1215),
.o01(east12_out1215),
.o02(west12_out1215),
.o03(north12_out1215),
.o04(south12_out1215)
);
router r13130
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in130),
.i01(east13_in130),
.i02(west13_in130),
.i03(north13_in130),
.i04(south13_in130),
.o00(local13_out130),
.o01(east13_out130),
.o02(west13_out130),
.o03(north13_out130),
.o04(south13_out130)
);
router r13131
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in131),
.i01(east13_in131),
.i02(west13_in131),
.i03(north13_in131),
.i04(south13_in131),
.o00(local13_out131),
.o01(east13_out131),
.o02(west13_out131),
.o03(north13_out131),
.o04(south13_out131)
);
router r13132
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in132),
.i01(east13_in132),
.i02(west13_in132),
.i03(north13_in132),
.i04(south13_in132),
.o00(local13_out132),
.o01(east13_out132),
.o02(west13_out132),
.o03(north13_out132),
.o04(south13_out132)
);
router r13133
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in133),
.i01(east13_in133),
.i02(west13_in133),
.i03(north13_in133),
.i04(south13_in133),
.o00(local13_out133),
.o01(east13_out133),
.o02(west13_out133),
.o03(north13_out133),
.o04(south13_out133)
);
router r13134
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in134),
.i01(east13_in134),
.i02(west13_in134),
.i03(north13_in134),
.i04(south13_in134),
.o00(local13_out134),
.o01(east13_out134),
.o02(west13_out134),
.o03(north13_out134),
.o04(south13_out134)
);
router r13135
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in135),
.i01(east13_in135),
.i02(west13_in135),
.i03(north13_in135),
.i04(south13_in135),
.o00(local13_out135),
.o01(east13_out135),
.o02(west13_out135),
.o03(north13_out135),
.o04(south13_out135)
);
router r13136
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in136),
.i01(east13_in136),
.i02(west13_in136),
.i03(north13_in136),
.i04(south13_in136),
.o00(local13_out136),
.o01(east13_out136),
.o02(west13_out136),
.o03(north13_out136),
.o04(south13_out136)
);
router r13137
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in137),
.i01(east13_in137),
.i02(west13_in137),
.i03(north13_in137),
.i04(south13_in137),
.o00(local13_out137),
.o01(east13_out137),
.o02(west13_out137),
.o03(north13_out137),
.o04(south13_out137)
);
router r13138
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in138),
.i01(east13_in138),
.i02(west13_in138),
.i03(north13_in138),
.i04(south13_in138),
.o00(local13_out138),
.o01(east13_out138),
.o02(west13_out138),
.o03(north13_out138),
.o04(south13_out138)
);
router r13139
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in139),
.i01(east13_in139),
.i02(west13_in139),
.i03(north13_in139),
.i04(south13_in139),
.o00(local13_out139),
.o01(east13_out139),
.o02(west13_out139),
.o03(north13_out139),
.o04(south13_out139)
);
router r131310
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in1310),
.i01(east13_in1310),
.i02(west13_in1310),
.i03(north13_in1310),
.i04(south13_in1310),
.o00(local13_out1310),
.o01(east13_out1310),
.o02(west13_out1310),
.o03(north13_out1310),
.o04(south13_out1310)
);
router r131311
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in1311),
.i01(east13_in1311),
.i02(west13_in1311),
.i03(north13_in1311),
.i04(south13_in1311),
.o00(local13_out1311),
.o01(east13_out1311),
.o02(west13_out1311),
.o03(north13_out1311),
.o04(south13_out1311)
);
router r131312
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in1312),
.i01(east13_in1312),
.i02(west13_in1312),
.i03(north13_in1312),
.i04(south13_in1312),
.o00(local13_out1312),
.o01(east13_out1312),
.o02(west13_out1312),
.o03(north13_out1312),
.o04(south13_out1312)
);
router r131313
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in1313),
.i01(east13_in1313),
.i02(west13_in1313),
.i03(north13_in1313),
.i04(south13_in1313),
.o00(local13_out1313),
.o01(east13_out1313),
.o02(west13_out1313),
.o03(north13_out1313),
.o04(south13_out1313)
);
router r131314
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in1314),
.i01(east13_in1314),
.i02(west13_in1314),
.i03(north13_in1314),
.i04(south13_in1314),
.o00(local13_out1314),
.o01(east13_out1314),
.o02(west13_out1314),
.o03(north13_out1314),
.o04(south13_out1314)
);
router r131315
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in1315),
.i01(east13_in1315),
.i02(west13_in1315),
.i03(north13_in1315),
.i04(south13_in1315),
.o00(local13_out1315),
.o01(east13_out1315),
.o02(west13_out1315),
.o03(north13_out1315),
.o04(south13_out1315)
);
router r14140
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in140),
.i01(east14_in140),
.i02(west14_in140),
.i03(north14_in140),
.i04(south14_in140),
.o00(local14_out140),
.o01(east14_out140),
.o02(west14_out140),
.o03(north14_out140),
.o04(south14_out140)
);
router r14141
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in141),
.i01(east14_in141),
.i02(west14_in141),
.i03(north14_in141),
.i04(south14_in141),
.o00(local14_out141),
.o01(east14_out141),
.o02(west14_out141),
.o03(north14_out141),
.o04(south14_out141)
);
router r14142
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in142),
.i01(east14_in142),
.i02(west14_in142),
.i03(north14_in142),
.i04(south14_in142),
.o00(local14_out142),
.o01(east14_out142),
.o02(west14_out142),
.o03(north14_out142),
.o04(south14_out142)
);
router r14143
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in143),
.i01(east14_in143),
.i02(west14_in143),
.i03(north14_in143),
.i04(south14_in143),
.o00(local14_out143),
.o01(east14_out143),
.o02(west14_out143),
.o03(north14_out143),
.o04(south14_out143)
);
router r14144
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in144),
.i01(east14_in144),
.i02(west14_in144),
.i03(north14_in144),
.i04(south14_in144),
.o00(local14_out144),
.o01(east14_out144),
.o02(west14_out144),
.o03(north14_out144),
.o04(south14_out144)
);
router r14145
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in145),
.i01(east14_in145),
.i02(west14_in145),
.i03(north14_in145),
.i04(south14_in145),
.o00(local14_out145),
.o01(east14_out145),
.o02(west14_out145),
.o03(north14_out145),
.o04(south14_out145)
);
router r14146
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in146),
.i01(east14_in146),
.i02(west14_in146),
.i03(north14_in146),
.i04(south14_in146),
.o00(local14_out146),
.o01(east14_out146),
.o02(west14_out146),
.o03(north14_out146),
.o04(south14_out146)
);
router r14147
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in147),
.i01(east14_in147),
.i02(west14_in147),
.i03(north14_in147),
.i04(south14_in147),
.o00(local14_out147),
.o01(east14_out147),
.o02(west14_out147),
.o03(north14_out147),
.o04(south14_out147)
);
router r14148
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in148),
.i01(east14_in148),
.i02(west14_in148),
.i03(north14_in148),
.i04(south14_in148),
.o00(local14_out148),
.o01(east14_out148),
.o02(west14_out148),
.o03(north14_out148),
.o04(south14_out148)
);
router r14149
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in149),
.i01(east14_in149),
.i02(west14_in149),
.i03(north14_in149),
.i04(south14_in149),
.o00(local14_out149),
.o01(east14_out149),
.o02(west14_out149),
.o03(north14_out149),
.o04(south14_out149)
);
router r141410
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in1410),
.i01(east14_in1410),
.i02(west14_in1410),
.i03(north14_in1410),
.i04(south14_in1410),
.o00(local14_out1410),
.o01(east14_out1410),
.o02(west14_out1410),
.o03(north14_out1410),
.o04(south14_out1410)
);
router r141411
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in1411),
.i01(east14_in1411),
.i02(west14_in1411),
.i03(north14_in1411),
.i04(south14_in1411),
.o00(local14_out1411),
.o01(east14_out1411),
.o02(west14_out1411),
.o03(north14_out1411),
.o04(south14_out1411)
);
router r141412
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in1412),
.i01(east14_in1412),
.i02(west14_in1412),
.i03(north14_in1412),
.i04(south14_in1412),
.o00(local14_out1412),
.o01(east14_out1412),
.o02(west14_out1412),
.o03(north14_out1412),
.o04(south14_out1412)
);
router r141413
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in1413),
.i01(east14_in1413),
.i02(west14_in1413),
.i03(north14_in1413),
.i04(south14_in1413),
.o00(local14_out1413),
.o01(east14_out1413),
.o02(west14_out1413),
.o03(north14_out1413),
.o04(south14_out1413)
);
router r141414
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in1414),
.i01(east14_in1414),
.i02(west14_in1414),
.i03(north14_in1414),
.i04(south14_in1414),
.o00(local14_out1414),
.o01(east14_out1414),
.o02(west14_out1414),
.o03(north14_out1414),
.o04(south14_out1414)
);
router r141415
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in1415),
.i01(east14_in1415),
.i02(west14_in1415),
.i03(north14_in1415),
.i04(south14_in1415),
.o00(local14_out1415),
.o01(east14_out1415),
.o02(west14_out1415),
.o03(north14_out1415),
.o04(south14_out1415)
);
router r15150
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in150),
.i01(east15_in150),
.i02(west15_in150),
.i03(north15_in150),
.i04(south15_in150),
.o00(local15_out150),
.o01(east15_out150),
.o02(west15_out150),
.o03(north15_out150),
.o04(south15_out150)
);
router r15151
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in151),
.i01(east15_in151),
.i02(west15_in151),
.i03(north15_in151),
.i04(south15_in151),
.o00(local15_out151),
.o01(east15_out151),
.o02(west15_out151),
.o03(north15_out151),
.o04(south15_out151)
);
router r15152
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in152),
.i01(east15_in152),
.i02(west15_in152),
.i03(north15_in152),
.i04(south15_in152),
.o00(local15_out152),
.o01(east15_out152),
.o02(west15_out152),
.o03(north15_out152),
.o04(south15_out152)
);
router r15153
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in153),
.i01(east15_in153),
.i02(west15_in153),
.i03(north15_in153),
.i04(south15_in153),
.o00(local15_out153),
.o01(east15_out153),
.o02(west15_out153),
.o03(north15_out153),
.o04(south15_out153)
);
router r15154
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in154),
.i01(east15_in154),
.i02(west15_in154),
.i03(north15_in154),
.i04(south15_in154),
.o00(local15_out154),
.o01(east15_out154),
.o02(west15_out154),
.o03(north15_out154),
.o04(south15_out154)
);
router r15155
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in155),
.i01(east15_in155),
.i02(west15_in155),
.i03(north15_in155),
.i04(south15_in155),
.o00(local15_out155),
.o01(east15_out155),
.o02(west15_out155),
.o03(north15_out155),
.o04(south15_out155)
);
router r15156
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in156),
.i01(east15_in156),
.i02(west15_in156),
.i03(north15_in156),
.i04(south15_in156),
.o00(local15_out156),
.o01(east15_out156),
.o02(west15_out156),
.o03(north15_out156),
.o04(south15_out156)
);
router r15157
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in157),
.i01(east15_in157),
.i02(west15_in157),
.i03(north15_in157),
.i04(south15_in157),
.o00(local15_out157),
.o01(east15_out157),
.o02(west15_out157),
.o03(north15_out157),
.o04(south15_out157)
);
router r15158
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in158),
.i01(east15_in158),
.i02(west15_in158),
.i03(north15_in158),
.i04(south15_in158),
.o00(local15_out158),
.o01(east15_out158),
.o02(west15_out158),
.o03(north15_out158),
.o04(south15_out158)
);
router r15159
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in159),
.i01(east15_in159),
.i02(west15_in159),
.i03(north15_in159),
.i04(south15_in159),
.o00(local15_out159),
.o01(east15_out159),
.o02(west15_out159),
.o03(north15_out159),
.o04(south15_out159)
);
router r151510
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in1510),
.i01(east15_in1510),
.i02(west15_in1510),
.i03(north15_in1510),
.i04(south15_in1510),
.o00(local15_out1510),
.o01(east15_out1510),
.o02(west15_out1510),
.o03(north15_out1510),
.o04(south15_out1510)
);
router r151511
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in1511),
.i01(east15_in1511),
.i02(west15_in1511),
.i03(north15_in1511),
.i04(south15_in1511),
.o00(local15_out1511),
.o01(east15_out1511),
.o02(west15_out1511),
.o03(north15_out1511),
.o04(south15_out1511)
);
router r151512
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in1512),
.i01(east15_in1512),
.i02(west15_in1512),
.i03(north15_in1512),
.i04(south15_in1512),
.o00(local15_out1512),
.o01(east15_out1512),
.o02(west15_out1512),
.o03(north15_out1512),
.o04(south15_out1512)
);
router r151513
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in1513),
.i01(east15_in1513),
.i02(west15_in1513),
.i03(north15_in1513),
.i04(south15_in1513),
.o00(local15_out1513),
.o01(east15_out1513),
.o02(west15_out1513),
.o03(north15_out1513),
.o04(south15_out1513)
);
router r151514
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in1514),
.i01(east15_in1514),
.i02(west15_in1514),
.i03(north15_in1514),
.i04(south15_in1514),
.o00(local15_out1514),
.o01(east15_out1514),
.o02(west15_out1514),
.o03(north15_out1514),
.o04(south15_out1514)
);
router r151515
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in1515),
.i01(east15_in1515),
.i02(west15_in1515),
.i03(north15_in1515),
.i04(south15_in1515),
.o00(local15_out1515),
.o01(east15_out1515),
.o02(west15_out1515),
.o03(north15_out1515),
.o04(south15_out1515)
);
always @ ( posedge clk)
begin
west0_in01<=east0_out00;
east0_in015<=west0_out00;
south15_in150<=north0_out00;
north1_in10<=south0_out00;
west0_in02<=east0_out01;
east0_in00<=west0_out01;
north1_in11<=south0_out01;
south15_in151<=north0_out01;
west0_in03<=east0_out02;
east0_in01<=west0_out02;
north1_in12<=south0_out02;
south15_in152<=north0_out02;
west0_in04<=east0_out03;
east0_in02<=west0_out03;
north1_in13<=south0_out03;
south15_in153<=north0_out03;
west0_in05<=east0_out04;
east0_in03<=west0_out04;
north1_in14<=south0_out04;
south15_in154<=north0_out04;
west0_in06<=east0_out05;
east0_in04<=west0_out05;
north1_in15<=south0_out05;
south15_in155<=north0_out05;
west0_in07<=east0_out06;
east0_in05<=west0_out06;
north1_in16<=south0_out06;
south15_in156<=north0_out06;
west0_in08<=east0_out07;
east0_in06<=west0_out07;
north1_in17<=south0_out07;
south15_in157<=north0_out07;
west0_in09<=east0_out08;
east0_in07<=west0_out08;
north1_in18<=south0_out08;
south15_in158<=north0_out08;
west0_in010<=east0_out09;
east0_in08<=west0_out09;
north1_in19<=south0_out09;
south15_in159<=north0_out09;
west0_in011<=east0_out010;
east0_in09<=west0_out010;
north1_in110<=south0_out010;
south15_in1510<=north0_out010;
west0_in012<=east0_out011;
east0_in010<=west0_out011;
north1_in111<=south0_out011;
south15_in1511<=north0_out011;
west0_in013<=east0_out012;
east0_in011<=west0_out012;
north1_in112<=south0_out012;
south15_in1512<=north0_out012;
west0_in014<=east0_out013;
east0_in012<=west0_out013;
north1_in113<=south0_out013;
south15_in1513<=north0_out013;
west0_in015<=east0_out014;
east0_in013<=west0_out014;
north1_in114<=south0_out014;
south15_in1514<=north0_out014;
west0_in00<=east0_out015;
east0_in014<=west0_out015;
north1_in115<=south0_out015;
south15_in1515<=north0_out015;
west1_in11<=east1_out10;
east1_in115<=west1_out10;
north2_in20<=south1_out10;
south0_in00<=north1_out10;
west1_in12<=east1_out11;
east1_in10<=west1_out11;
south0_in01<=north1_out11;
north2_in21<=south1_out11;
west1_in13<=east1_out12;
east1_in11<=west1_out12;
south0_in02<=north1_out12;
north2_in22<=south1_out12;
west1_in14<=east1_out13;
east1_in12<=west1_out13;
south0_in03<=north1_out13;
north2_in23<=south1_out13;
west1_in15<=east1_out14;
east1_in13<=west1_out14;
south0_in04<=north1_out14;
north2_in24<=south1_out14;
west1_in16<=east1_out15;
east1_in14<=west1_out15;
south0_in05<=north1_out15;
north2_in25<=south1_out15;
west1_in17<=east1_out16;
east1_in15<=west1_out16;
south0_in06<=north1_out16;
north2_in26<=south1_out16;
west1_in18<=east1_out17;
east1_in16<=west1_out17;
south0_in07<=north1_out17;
north2_in27<=south1_out17;
west1_in19<=east1_out18;
east1_in17<=west1_out18;
south0_in08<=north1_out18;
north2_in28<=south1_out18;
west1_in110<=east1_out19;
east1_in18<=west1_out19;
south0_in09<=north1_out19;
north2_in29<=south1_out19;
west1_in111<=east1_out110;
east1_in19<=west1_out110;
south0_in010<=north1_out110;
north2_in210<=south1_out110;
west1_in112<=east1_out111;
east1_in110<=west1_out111;
south0_in011<=north1_out111;
north2_in211<=south1_out111;
west1_in113<=east1_out112;
east1_in111<=west1_out112;
south0_in012<=north1_out112;
north2_in212<=south1_out112;
west1_in114<=east1_out113;
east1_in112<=west1_out113;
south0_in013<=north1_out113;
north2_in213<=south1_out113;
west1_in115<=east1_out114;
east1_in113<=west1_out114;
south0_in014<=north1_out114;
north2_in214<=south1_out114;
west1_in10<=east1_out115;
east1_in114<=west1_out115;
north2_in215<=south1_out115;
south0_in015<=north1_out115;
west2_in21<=east2_out20;
east2_in215<=west2_out20;
north3_in30<=south2_out20;
south1_in10<=north2_out20;
west2_in22<=east2_out21;
east2_in20<=west2_out21;
south1_in11<=north2_out21;
north3_in31<=south2_out21;
west2_in23<=east2_out22;
east2_in21<=west2_out22;
south1_in12<=north2_out22;
north3_in32<=south2_out22;
west2_in24<=east2_out23;
east2_in22<=west2_out23;
south1_in13<=north2_out23;
north3_in33<=south2_out23;
west2_in25<=east2_out24;
east2_in23<=west2_out24;
south1_in14<=north2_out24;
north3_in34<=south2_out24;
west2_in26<=east2_out25;
east2_in24<=west2_out25;
south1_in15<=north2_out25;
north3_in35<=south2_out25;
west2_in27<=east2_out26;
east2_in25<=west2_out26;
south1_in16<=north2_out26;
north3_in36<=south2_out26;
west2_in28<=east2_out27;
east2_in26<=west2_out27;
south1_in17<=north2_out27;
north3_in37<=south2_out27;
west2_in29<=east2_out28;
east2_in27<=west2_out28;
south1_in18<=north2_out28;
north3_in38<=south2_out28;
west2_in210<=east2_out29;
east2_in28<=west2_out29;
south1_in19<=north2_out29;
north3_in39<=south2_out29;
west2_in211<=east2_out210;
east2_in29<=west2_out210;
south1_in110<=north2_out210;
north3_in310<=south2_out210;
west2_in212<=east2_out211;
east2_in210<=west2_out211;
south1_in111<=north2_out211;
north3_in311<=south2_out211;
west2_in213<=east2_out212;
east2_in211<=west2_out212;
south1_in112<=north2_out212;
north3_in312<=south2_out212;
west2_in214<=east2_out213;
east2_in212<=west2_out213;
south1_in113<=north2_out213;
north3_in313<=south2_out213;
west2_in215<=east2_out214;
east2_in213<=west2_out214;
south1_in114<=north2_out214;
north3_in314<=south2_out214;
west2_in20<=east2_out215;
east2_in214<=west2_out215;
north3_in315<=south2_out215;
south1_in115<=north2_out215;
west3_in31<=east3_out30;
east3_in315<=west3_out30;
north4_in40<=south3_out30;
south2_in20<=north3_out30;
west3_in32<=east3_out31;
east3_in30<=west3_out31;
south2_in21<=north3_out31;
north4_in41<=south3_out31;
west3_in33<=east3_out32;
east3_in31<=west3_out32;
south2_in22<=north3_out32;
north4_in42<=south3_out32;
west3_in34<=east3_out33;
east3_in32<=west3_out33;
south2_in23<=north3_out33;
north4_in43<=south3_out33;
west3_in35<=east3_out34;
east3_in33<=west3_out34;
south2_in24<=north3_out34;
north4_in44<=south3_out34;
west3_in36<=east3_out35;
east3_in34<=west3_out35;
south2_in25<=north3_out35;
north4_in45<=south3_out35;
west3_in37<=east3_out36;
east3_in35<=west3_out36;
south2_in26<=north3_out36;
north4_in46<=south3_out36;
west3_in38<=east3_out37;
east3_in36<=west3_out37;
south2_in27<=north3_out37;
north4_in47<=south3_out37;
west3_in39<=east3_out38;
east3_in37<=west3_out38;
south2_in28<=north3_out38;
north4_in48<=south3_out38;
west3_in310<=east3_out39;
east3_in38<=west3_out39;
south2_in29<=north3_out39;
north4_in49<=south3_out39;
west3_in311<=east3_out310;
east3_in39<=west3_out310;
south2_in210<=north3_out310;
north4_in410<=south3_out310;
west3_in312<=east3_out311;
east3_in310<=west3_out311;
south2_in211<=north3_out311;
north4_in411<=south3_out311;
west3_in313<=east3_out312;
east3_in311<=west3_out312;
south2_in212<=north3_out312;
north4_in412<=south3_out312;
west3_in314<=east3_out313;
east3_in312<=west3_out313;
south2_in213<=north3_out313;
north4_in413<=south3_out313;
west3_in315<=east3_out314;
east3_in313<=west3_out314;
south2_in214<=north3_out314;
north4_in414<=south3_out314;
west3_in30<=east3_out315;
east3_in314<=west3_out315;
north4_in415<=south3_out315;
south2_in215<=north3_out315;
west4_in41<=east4_out40;
east4_in415<=west4_out40;
north5_in50<=south4_out40;
south3_in30<=north4_out40;
west4_in42<=east4_out41;
east4_in40<=west4_out41;
south3_in31<=north4_out41;
north5_in51<=south4_out41;
west4_in43<=east4_out42;
east4_in41<=west4_out42;
south3_in32<=north4_out42;
north5_in52<=south4_out42;
west4_in44<=east4_out43;
east4_in42<=west4_out43;
south3_in33<=north4_out43;
north5_in53<=south4_out43;
west4_in45<=east4_out44;
east4_in43<=west4_out44;
south3_in34<=north4_out44;
north5_in54<=south4_out44;
west4_in46<=east4_out45;
east4_in44<=west4_out45;
south3_in35<=north4_out45;
north5_in55<=south4_out45;
west4_in47<=east4_out46;
east4_in45<=west4_out46;
south3_in36<=north4_out46;
north5_in56<=south4_out46;
west4_in48<=east4_out47;
east4_in46<=west4_out47;
south3_in37<=north4_out47;
north5_in57<=south4_out47;
west4_in49<=east4_out48;
east4_in47<=west4_out48;
south3_in38<=north4_out48;
north5_in58<=south4_out48;
west4_in410<=east4_out49;
east4_in48<=west4_out49;
south3_in39<=north4_out49;
north5_in59<=south4_out49;
west4_in411<=east4_out410;
east4_in49<=west4_out410;
south3_in310<=north4_out410;
north5_in510<=south4_out410;
west4_in412<=east4_out411;
east4_in410<=west4_out411;
south3_in311<=north4_out411;
north5_in511<=south4_out411;
west4_in413<=east4_out412;
east4_in411<=west4_out412;
south3_in312<=north4_out412;
north5_in512<=south4_out412;
west4_in414<=east4_out413;
east4_in412<=west4_out413;
south3_in313<=north4_out413;
north5_in513<=south4_out413;
west4_in415<=east4_out414;
east4_in413<=west4_out414;
south3_in314<=north4_out414;
north5_in514<=south4_out414;
west4_in40<=east4_out415;
east4_in414<=west4_out415;
north5_in515<=south4_out415;
south3_in315<=north4_out415;
west5_in51<=east5_out50;
east5_in515<=west5_out50;
north6_in60<=south5_out50;
south4_in40<=north5_out50;
west5_in52<=east5_out51;
east5_in50<=west5_out51;
south4_in41<=north5_out51;
north6_in61<=south5_out51;
west5_in53<=east5_out52;
east5_in51<=west5_out52;
south4_in42<=north5_out52;
north6_in62<=south5_out52;
west5_in54<=east5_out53;
east5_in52<=west5_out53;
south4_in43<=north5_out53;
north6_in63<=south5_out53;
west5_in55<=east5_out54;
east5_in53<=west5_out54;
south4_in44<=north5_out54;
north6_in64<=south5_out54;
west5_in56<=east5_out55;
east5_in54<=west5_out55;
south4_in45<=north5_out55;
north6_in65<=south5_out55;
west5_in57<=east5_out56;
east5_in55<=west5_out56;
south4_in46<=north5_out56;
north6_in66<=south5_out56;
west5_in58<=east5_out57;
east5_in56<=west5_out57;
south4_in47<=north5_out57;
north6_in67<=south5_out57;
west5_in59<=east5_out58;
east5_in57<=west5_out58;
south4_in48<=north5_out58;
north6_in68<=south5_out58;
west5_in510<=east5_out59;
east5_in58<=west5_out59;
south4_in49<=north5_out59;
north6_in69<=south5_out59;
west5_in511<=east5_out510;
east5_in59<=west5_out510;
south4_in410<=north5_out510;
north6_in610<=south5_out510;
west5_in512<=east5_out511;
east5_in510<=west5_out511;
south4_in411<=north5_out511;
north6_in611<=south5_out511;
west5_in513<=east5_out512;
east5_in511<=west5_out512;
south4_in412<=north5_out512;
north6_in612<=south5_out512;
west5_in514<=east5_out513;
east5_in512<=west5_out513;
south4_in413<=north5_out513;
north6_in613<=south5_out513;
west5_in515<=east5_out514;
east5_in513<=west5_out514;
south4_in414<=north5_out514;
north6_in614<=south5_out514;
west5_in50<=east5_out515;
east5_in514<=west5_out515;
north6_in615<=south5_out515;
south4_in415<=north5_out515;
west6_in61<=east6_out60;
east6_in615<=west6_out60;
north7_in70<=south6_out60;
south5_in50<=north6_out60;
west6_in62<=east6_out61;
east6_in60<=west6_out61;
south5_in51<=north6_out61;
north7_in71<=south6_out61;
west6_in63<=east6_out62;
east6_in61<=west6_out62;
south5_in52<=north6_out62;
north7_in72<=south6_out62;
west6_in64<=east6_out63;
east6_in62<=west6_out63;
south5_in53<=north6_out63;
north7_in73<=south6_out63;
west6_in65<=east6_out64;
east6_in63<=west6_out64;
south5_in54<=north6_out64;
north7_in74<=south6_out64;
west6_in66<=east6_out65;
east6_in64<=west6_out65;
south5_in55<=north6_out65;
north7_in75<=south6_out65;
west6_in67<=east6_out66;
east6_in65<=west6_out66;
south5_in56<=north6_out66;
north7_in76<=south6_out66;
west6_in68<=east6_out67;
east6_in66<=west6_out67;
south5_in57<=north6_out67;
north7_in77<=south6_out67;
west6_in69<=east6_out68;
east6_in67<=west6_out68;
south5_in58<=north6_out68;
north7_in78<=south6_out68;
west6_in610<=east6_out69;
east6_in68<=west6_out69;
south5_in59<=north6_out69;
north7_in79<=south6_out69;
west6_in611<=east6_out610;
east6_in69<=west6_out610;
south5_in510<=north6_out610;
north7_in710<=south6_out610;
west6_in612<=east6_out611;
east6_in610<=west6_out611;
south5_in511<=north6_out611;
north7_in711<=south6_out611;
west6_in613<=east6_out612;
east6_in611<=west6_out612;
south5_in512<=north6_out612;
north7_in712<=south6_out612;
west6_in614<=east6_out613;
east6_in612<=west6_out613;
south5_in513<=north6_out613;
north7_in713<=south6_out613;
west6_in615<=east6_out614;
east6_in613<=west6_out614;
south5_in514<=north6_out614;
north7_in714<=south6_out614;
west6_in60<=east6_out615;
east6_in614<=west6_out615;
north7_in715<=south6_out615;
south5_in515<=north6_out615;
west7_in71<=east7_out70;
east7_in715<=west7_out70;
north8_in80<=south7_out70;
south6_in60<=north7_out70;
west7_in72<=east7_out71;
east7_in70<=west7_out71;
south6_in61<=north7_out71;
north8_in81<=south7_out71;
west7_in73<=east7_out72;
east7_in71<=west7_out72;
south6_in62<=north7_out72;
north8_in82<=south7_out72;
west7_in74<=east7_out73;
east7_in72<=west7_out73;
south6_in63<=north7_out73;
north8_in83<=south7_out73;
west7_in75<=east7_out74;
east7_in73<=west7_out74;
south6_in64<=north7_out74;
north8_in84<=south7_out74;
west7_in76<=east7_out75;
east7_in74<=west7_out75;
south6_in65<=north7_out75;
north8_in85<=south7_out75;
west7_in77<=east7_out76;
east7_in75<=west7_out76;
south6_in66<=north7_out76;
north8_in86<=south7_out76;
west7_in78<=east7_out77;
east7_in76<=west7_out77;
south6_in67<=north7_out77;
north8_in87<=south7_out77;
west7_in79<=east7_out78;
east7_in77<=west7_out78;
south6_in68<=north7_out78;
north8_in88<=south7_out78;
west7_in710<=east7_out79;
east7_in78<=west7_out79;
south6_in69<=north7_out79;
north8_in89<=south7_out79;
west7_in711<=east7_out710;
east7_in79<=west7_out710;
south6_in610<=north7_out710;
north8_in810<=south7_out710;
west7_in712<=east7_out711;
east7_in710<=west7_out711;
south6_in611<=north7_out711;
north8_in811<=south7_out711;
west7_in713<=east7_out712;
east7_in711<=west7_out712;
south6_in612<=north7_out712;
north8_in812<=south7_out712;
west7_in714<=east7_out713;
east7_in712<=west7_out713;
south6_in613<=north7_out713;
north8_in813<=south7_out713;
west7_in715<=east7_out714;
east7_in713<=west7_out714;
south6_in614<=north7_out714;
north8_in814<=south7_out714;
west7_in70<=east7_out715;
east7_in714<=west7_out715;
north8_in815<=south7_out715;
south6_in615<=north7_out715;
west8_in81<=east8_out80;
east8_in815<=west8_out80;
north9_in90<=south8_out80;
south7_in70<=north8_out80;
west8_in82<=east8_out81;
east8_in80<=west8_out81;
south7_in71<=north8_out81;
north9_in91<=south8_out81;
west8_in83<=east8_out82;
east8_in81<=west8_out82;
south7_in72<=north8_out82;
north9_in92<=south8_out82;
west8_in84<=east8_out83;
east8_in82<=west8_out83;
south7_in73<=north8_out83;
north9_in93<=south8_out83;
west8_in85<=east8_out84;
east8_in83<=west8_out84;
south7_in74<=north8_out84;
north9_in94<=south8_out84;
west8_in86<=east8_out85;
east8_in84<=west8_out85;
south7_in75<=north8_out85;
north9_in95<=south8_out85;
west8_in87<=east8_out86;
east8_in85<=west8_out86;
south7_in76<=north8_out86;
north9_in96<=south8_out86;
west8_in88<=east8_out87;
east8_in86<=west8_out87;
south7_in77<=north8_out87;
north9_in97<=south8_out87;
west8_in89<=east8_out88;
east8_in87<=west8_out88;
south7_in78<=north8_out88;
north9_in98<=south8_out88;
west8_in810<=east8_out89;
east8_in88<=west8_out89;
south7_in79<=north8_out89;
north9_in99<=south8_out89;
west8_in811<=east8_out810;
east8_in89<=west8_out810;
south7_in710<=north8_out810;
north9_in910<=south8_out810;
west8_in812<=east8_out811;
east8_in810<=west8_out811;
south7_in711<=north8_out811;
north9_in911<=south8_out811;
west8_in813<=east8_out812;
east8_in811<=west8_out812;
south7_in712<=north8_out812;
north9_in912<=south8_out812;
west8_in814<=east8_out813;
east8_in812<=west8_out813;
south7_in713<=north8_out813;
north9_in913<=south8_out813;
west8_in815<=east8_out814;
east8_in813<=west8_out814;
south7_in714<=north8_out814;
north9_in914<=south8_out814;
west8_in80<=east8_out815;
east8_in814<=west8_out815;
north9_in915<=south8_out815;
south7_in715<=north8_out815;
west9_in91<=east9_out90;
east9_in915<=west9_out90;
north10_in100<=south9_out90;
south8_in80<=north9_out90;
west9_in92<=east9_out91;
east9_in90<=west9_out91;
south8_in81<=north9_out91;
north10_in101<=south9_out91;
west9_in93<=east9_out92;
east9_in91<=west9_out92;
south8_in82<=north9_out92;
north10_in102<=south9_out92;
west9_in94<=east9_out93;
east9_in92<=west9_out93;
south8_in83<=north9_out93;
north10_in103<=south9_out93;
west9_in95<=east9_out94;
east9_in93<=west9_out94;
south8_in84<=north9_out94;
north10_in104<=south9_out94;
west9_in96<=east9_out95;
east9_in94<=west9_out95;
south8_in85<=north9_out95;
north10_in105<=south9_out95;
west9_in97<=east9_out96;
east9_in95<=west9_out96;
south8_in86<=north9_out96;
north10_in106<=south9_out96;
west9_in98<=east9_out97;
east9_in96<=west9_out97;
south8_in87<=north9_out97;
north10_in107<=south9_out97;
west9_in99<=east9_out98;
east9_in97<=west9_out98;
south8_in88<=north9_out98;
north10_in108<=south9_out98;
west9_in910<=east9_out99;
east9_in98<=west9_out99;
south8_in89<=north9_out99;
north10_in109<=south9_out99;
west9_in911<=east9_out910;
east9_in99<=west9_out910;
south8_in810<=north9_out910;
north10_in1010<=south9_out910;
west9_in912<=east9_out911;
east9_in910<=west9_out911;
south8_in811<=north9_out911;
north10_in1011<=south9_out911;
west9_in913<=east9_out912;
east9_in911<=west9_out912;
south8_in812<=north9_out912;
north10_in1012<=south9_out912;
west9_in914<=east9_out913;
east9_in912<=west9_out913;
south8_in813<=north9_out913;
north10_in1013<=south9_out913;
west9_in915<=east9_out914;
east9_in913<=west9_out914;
south8_in814<=north9_out914;
north10_in1014<=south9_out914;
west9_in90<=east9_out915;
east9_in914<=west9_out915;
north10_in1015<=south9_out915;
south8_in815<=north9_out915;
west10_in101<=east10_out100;
east10_in1015<=west10_out100;
north11_in110<=south10_out100;
south9_in90<=north10_out100;
west10_in102<=east10_out101;
east10_in100<=west10_out101;
south9_in91<=north10_out101;
north11_in111<=south10_out101;
west10_in103<=east10_out102;
east10_in101<=west10_out102;
south9_in92<=north10_out102;
north11_in112<=south10_out102;
west10_in104<=east10_out103;
east10_in102<=west10_out103;
south9_in93<=north10_out103;
north11_in113<=south10_out103;
west10_in105<=east10_out104;
east10_in103<=west10_out104;
south9_in94<=north10_out104;
north11_in114<=south10_out104;
west10_in106<=east10_out105;
east10_in104<=west10_out105;
south9_in95<=north10_out105;
north11_in115<=south10_out105;
west10_in107<=east10_out106;
east10_in105<=west10_out106;
south9_in96<=north10_out106;
north11_in116<=south10_out106;
west10_in108<=east10_out107;
east10_in106<=west10_out107;
south9_in97<=north10_out107;
north11_in117<=south10_out107;
west10_in109<=east10_out108;
east10_in107<=west10_out108;
south9_in98<=north10_out108;
north11_in118<=south10_out108;
west10_in1010<=east10_out109;
east10_in108<=west10_out109;
south9_in99<=north10_out109;
north11_in119<=south10_out109;
west10_in1011<=east10_out1010;
east10_in109<=west10_out1010;
south9_in910<=north10_out1010;
north11_in1110<=south10_out1010;
west10_in1012<=east10_out1011;
east10_in1010<=west10_out1011;
south9_in911<=north10_out1011;
north11_in1111<=south10_out1011;
west10_in1013<=east10_out1012;
east10_in1011<=west10_out1012;
south9_in912<=north10_out1012;
north11_in1112<=south10_out1012;
west10_in1014<=east10_out1013;
east10_in1012<=west10_out1013;
south9_in913<=north10_out1013;
north11_in1113<=south10_out1013;
west10_in1015<=east10_out1014;
east10_in1013<=west10_out1014;
south9_in914<=north10_out1014;
north11_in1114<=south10_out1014;
west10_in100<=east10_out1015;
east10_in1014<=west10_out1015;
north11_in1115<=south10_out1015;
south9_in915<=north10_out1015;
west11_in111<=east11_out110;
east11_in1115<=west11_out110;
north12_in120<=south11_out110;
south10_in100<=north11_out110;
west11_in112<=east11_out111;
east11_in110<=west11_out111;
south10_in101<=north11_out111;
north12_in121<=south11_out111;
west11_in113<=east11_out112;
east11_in111<=west11_out112;
south10_in102<=north11_out112;
north12_in122<=south11_out112;
west11_in114<=east11_out113;
east11_in112<=west11_out113;
south10_in103<=north11_out113;
north12_in123<=south11_out113;
west11_in115<=east11_out114;
east11_in113<=west11_out114;
south10_in104<=north11_out114;
north12_in124<=south11_out114;
west11_in116<=east11_out115;
east11_in114<=west11_out115;
south10_in105<=north11_out115;
north12_in125<=south11_out115;
west11_in117<=east11_out116;
east11_in115<=west11_out116;
south10_in106<=north11_out116;
north12_in126<=south11_out116;
west11_in118<=east11_out117;
east11_in116<=west11_out117;
south10_in107<=north11_out117;
north12_in127<=south11_out117;
west11_in119<=east11_out118;
east11_in117<=west11_out118;
south10_in108<=north11_out118;
north12_in128<=south11_out118;
west11_in1110<=east11_out119;
east11_in118<=west11_out119;
south10_in109<=north11_out119;
north12_in129<=south11_out119;
west11_in1111<=east11_out1110;
east11_in119<=west11_out1110;
south10_in1010<=north11_out1110;
north12_in1210<=south11_out1110;
west11_in1112<=east11_out1111;
east11_in1110<=west11_out1111;
south10_in1011<=north11_out1111;
north12_in1211<=south11_out1111;
west11_in1113<=east11_out1112;
east11_in1111<=west11_out1112;
south10_in1012<=north11_out1112;
north12_in1212<=south11_out1112;
west11_in1114<=east11_out1113;
east11_in1112<=west11_out1113;
south10_in1013<=north11_out1113;
north12_in1213<=south11_out1113;
west11_in1115<=east11_out1114;
east11_in1113<=west11_out1114;
south10_in1014<=north11_out1114;
north12_in1214<=south11_out1114;
west11_in110<=east11_out1115;
east11_in1114<=west11_out1115;
north12_in1215<=south11_out1115;
south10_in1015<=north11_out1115;
west12_in121<=east12_out120;
east12_in1215<=west12_out120;
north13_in130<=south12_out120;
south11_in110<=north12_out120;
west12_in122<=east12_out121;
east12_in120<=west12_out121;
south11_in111<=north12_out121;
north13_in131<=south12_out121;
west12_in123<=east12_out122;
east12_in121<=west12_out122;
south11_in112<=north12_out122;
north13_in132<=south12_out122;
west12_in124<=east12_out123;
east12_in122<=west12_out123;
south11_in113<=north12_out123;
north13_in133<=south12_out123;
west12_in125<=east12_out124;
east12_in123<=west12_out124;
south11_in114<=north12_out124;
north13_in134<=south12_out124;
west12_in126<=east12_out125;
east12_in124<=west12_out125;
south11_in115<=north12_out125;
north13_in135<=south12_out125;
west12_in127<=east12_out126;
east12_in125<=west12_out126;
south11_in116<=north12_out126;
north13_in136<=south12_out126;
west12_in128<=east12_out127;
east12_in126<=west12_out127;
south11_in117<=north12_out127;
north13_in137<=south12_out127;
west12_in129<=east12_out128;
east12_in127<=west12_out128;
south11_in118<=north12_out128;
north13_in138<=south12_out128;
west12_in1210<=east12_out129;
east12_in128<=west12_out129;
south11_in119<=north12_out129;
north13_in139<=south12_out129;
west12_in1211<=east12_out1210;
east12_in129<=west12_out1210;
south11_in1110<=north12_out1210;
north13_in1310<=south12_out1210;
west12_in1212<=east12_out1211;
east12_in1210<=west12_out1211;
south11_in1111<=north12_out1211;
north13_in1311<=south12_out1211;
west12_in1213<=east12_out1212;
east12_in1211<=west12_out1212;
south11_in1112<=north12_out1212;
north13_in1312<=south12_out1212;
west12_in1214<=east12_out1213;
east12_in1212<=west12_out1213;
south11_in1113<=north12_out1213;
north13_in1313<=south12_out1213;
west12_in1215<=east12_out1214;
east12_in1213<=west12_out1214;
south11_in1114<=north12_out1214;
north13_in1314<=south12_out1214;
west12_in120<=east12_out1215;
east12_in1214<=west12_out1215;
north13_in1315<=south12_out1215;
south11_in1115<=north12_out1215;
west13_in131<=east13_out130;
east13_in1315<=west13_out130;
north14_in140<=south13_out130;
south12_in120<=north13_out130;
west13_in132<=east13_out131;
east13_in130<=west13_out131;
south12_in121<=north13_out131;
north14_in141<=south13_out131;
west13_in133<=east13_out132;
east13_in131<=west13_out132;
south12_in122<=north13_out132;
north14_in142<=south13_out132;
west13_in134<=east13_out133;
east13_in132<=west13_out133;
south12_in123<=north13_out133;
north14_in143<=south13_out133;
west13_in135<=east13_out134;
east13_in133<=west13_out134;
south12_in124<=north13_out134;
north14_in144<=south13_out134;
west13_in136<=east13_out135;
east13_in134<=west13_out135;
south12_in125<=north13_out135;
north14_in145<=south13_out135;
west13_in137<=east13_out136;
east13_in135<=west13_out136;
south12_in126<=north13_out136;
north14_in146<=south13_out136;
west13_in138<=east13_out137;
east13_in136<=west13_out137;
south12_in127<=north13_out137;
north14_in147<=south13_out137;
west13_in139<=east13_out138;
east13_in137<=west13_out138;
south12_in128<=north13_out138;
north14_in148<=south13_out138;
west13_in1310<=east13_out139;
east13_in138<=west13_out139;
south12_in129<=north13_out139;
north14_in149<=south13_out139;
west13_in1311<=east13_out1310;
east13_in139<=west13_out1310;
south12_in1210<=north13_out1310;
north14_in1410<=south13_out1310;
west13_in1312<=east13_out1311;
east13_in1310<=west13_out1311;
south12_in1211<=north13_out1311;
north14_in1411<=south13_out1311;
west13_in1313<=east13_out1312;
east13_in1311<=west13_out1312;
south12_in1212<=north13_out1312;
north14_in1412<=south13_out1312;
west13_in1314<=east13_out1313;
east13_in1312<=west13_out1313;
south12_in1213<=north13_out1313;
north14_in1413<=south13_out1313;
west13_in1315<=east13_out1314;
east13_in1313<=west13_out1314;
south12_in1214<=north13_out1314;
north14_in1414<=south13_out1314;
west13_in130<=east13_out1315;
east13_in1314<=west13_out1315;
north14_in1415<=south13_out1315;
south12_in1215<=north13_out1315;
west14_in141<=east14_out140;
east14_in1415<=west14_out140;
north15_in150<=south14_out140;
south13_in130<=north14_out140;
west14_in142<=east14_out141;
east14_in140<=west14_out141;
south13_in131<=north14_out141;
north15_in151<=south14_out141;
west14_in143<=east14_out142;
east14_in141<=west14_out142;
south13_in132<=north14_out142;
north15_in152<=south14_out142;
west14_in144<=east14_out143;
east14_in142<=west14_out143;
south13_in133<=north14_out143;
north15_in153<=south14_out143;
west14_in145<=east14_out144;
east14_in143<=west14_out144;
south13_in134<=north14_out144;
north15_in154<=south14_out144;
west14_in146<=east14_out145;
east14_in144<=west14_out145;
south13_in135<=north14_out145;
north15_in155<=south14_out145;
west14_in147<=east14_out146;
east14_in145<=west14_out146;
south13_in136<=north14_out146;
north15_in156<=south14_out146;
west14_in148<=east14_out147;
east14_in146<=west14_out147;
south13_in137<=north14_out147;
north15_in157<=south14_out147;
west14_in149<=east14_out148;
east14_in147<=west14_out148;
south13_in138<=north14_out148;
north15_in158<=south14_out148;
west14_in1410<=east14_out149;
east14_in148<=west14_out149;
south13_in139<=north14_out149;
north15_in159<=south14_out149;
west14_in1411<=east14_out1410;
east14_in149<=west14_out1410;
south13_in1310<=north14_out1410;
north15_in1510<=south14_out1410;
west14_in1412<=east14_out1411;
east14_in1410<=west14_out1411;
south13_in1311<=north14_out1411;
north15_in1511<=south14_out1411;
west14_in1413<=east14_out1412;
east14_in1411<=west14_out1412;
south13_in1312<=north14_out1412;
north15_in1512<=south14_out1412;
west14_in1414<=east14_out1413;
east14_in1412<=west14_out1413;
south13_in1313<=north14_out1413;
north15_in1513<=south14_out1413;
west14_in1415<=east14_out1414;
east14_in1413<=west14_out1414;
south13_in1314<=north14_out1414;
north15_in1514<=south14_out1414;
west14_in140<=east14_out1415;
east14_in1414<=west14_out1415;
north15_in1515<=south14_out1415;
south13_in1315<=north14_out1415;
west15_in151<=east15_out150;
east15_in1515<=west15_out150;
north0_in00<=south15_out150;
south14_in140<=north15_out150;
west15_in152<=east15_out151;
east15_in150<=west15_out151;
south0_in01<=south15_out151;
south14_in141<=north15_out151;
west15_in153<=east15_out152;
east15_in151<=west15_out152;
south0_in02<=south15_out152;
south14_in142<=north15_out152;
west15_in154<=east15_out153;
east15_in152<=west15_out153;
south0_in03<=south15_out153;
south14_in143<=north15_out153;
west15_in155<=east15_out154;
east15_in153<=west15_out154;
south0_in04<=south15_out154;
south14_in144<=north15_out154;
west15_in156<=east15_out155;
east15_in154<=west15_out155;
south0_in05<=south15_out155;
south14_in145<=north15_out155;
west15_in157<=east15_out156;
east15_in155<=west15_out156;
south0_in06<=south15_out156;
south14_in146<=north15_out156;
west15_in158<=east15_out157;
east15_in156<=west15_out157;
south0_in07<=south15_out157;
south14_in147<=north15_out157;
west15_in159<=east15_out158;
east15_in157<=west15_out158;
south0_in08<=south15_out158;
south14_in148<=north15_out158;
west15_in1510<=east15_out159;
east15_in158<=west15_out159;
south0_in09<=south15_out159;
south14_in149<=north15_out159;
west15_in1511<=east15_out1510;
east15_in159<=west15_out1510;
south0_in010<=south15_out1510;
south14_in1410<=north15_out1510;
west15_in1512<=east15_out1511;
east15_in1510<=west15_out1511;
south0_in011<=south15_out1511;
south14_in1411<=north15_out1511;
west15_in1513<=east15_out1512;
east15_in1511<=west15_out1512;
south0_in012<=south15_out1512;
south14_in1412<=north15_out1512;
west15_in1514<=east15_out1513;
east15_in1512<=west15_out1513;
south0_in013<=south15_out1513;
south14_in1413<=north15_out1513;
west15_in1515<=east15_out1514;
east15_in1513<=west15_out1514;
south0_in014<=south15_out1514;
south14_in1414<=north15_out1514;
west15_in150<=east15_out1515;
east15_in1514<=west15_out1515;
north0_in015<=south15_out1515;
south14_in1415<=north15_out1515;
end
endmodule
