module test_case_1 #(parameter NUM_AGENT=6,
                               PIPE_DLY =4,
                               N = 10,
                               M = 20
                    ) 
                       (
                            randomignore
                            input                   [0:2]     clk [10:8];
                            input                             rst_n
                            input  logic [NUM_AGENT-1:0] req,
                            output logic [NUM_AGENT-1:0] gnt,
                            output logic [2:0]           arbiter_state,
                            output                       arb_idle,
                                                         arb_busy
                            abc.xyz [2:0] shabalaba
                       ) ;
bla bla
bla bla
bla bla
bla bla
bla bla
bla bla
bla bla
bla bla
bla bla
bla bla

endmodule

