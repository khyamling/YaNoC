module torus (
local0_in00,local0_out00,
local0_in01,local0_out01,
local0_in02,local0_out02,
local0_in03,local0_out03,
local0_in04,local0_out04,
local0_in05,local0_out05,
local0_in06,local0_out06,
local0_in07,local0_out07,
local0_in08,local0_out08,
local0_in09,local0_out09,
local1_in10,local1_out10,
local1_in11,local1_out11,
local1_in12,local1_out12,
local1_in13,local1_out13,
local1_in14,local1_out14,
local1_in15,local1_out15,
local1_in16,local1_out16,
local1_in17,local1_out17,
local1_in18,local1_out18,
local1_in19,local1_out19,
local2_in20,local2_out20,
local2_in21,local2_out21,
local2_in22,local2_out22,
local2_in23,local2_out23,
local2_in24,local2_out24,
local2_in25,local2_out25,
local2_in26,local2_out26,
local2_in27,local2_out27,
local2_in28,local2_out28,
local2_in29,local2_out29,
local3_in30,local3_out30,
local3_in31,local3_out31,
local3_in32,local3_out32,
local3_in33,local3_out33,
local3_in34,local3_out34,
local3_in35,local3_out35,
local3_in36,local3_out36,
local3_in37,local3_out37,
local3_in38,local3_out38,
local3_in39,local3_out39,
local4_in40,local4_out40,
local4_in41,local4_out41,
local4_in42,local4_out42,
local4_in43,local4_out43,
local4_in44,local4_out44,
local4_in45,local4_out45,
local4_in46,local4_out46,
local4_in47,local4_out47,
local4_in48,local4_out48,
local4_in49,local4_out49,
local5_in50,local5_out50,
local5_in51,local5_out51,
local5_in52,local5_out52,
local5_in53,local5_out53,
local5_in54,local5_out54,
local5_in55,local5_out55,
local5_in56,local5_out56,
local5_in57,local5_out57,
local5_in58,local5_out58,
local5_in59,local5_out59,
local6_in60,local6_out60,
local6_in61,local6_out61,
local6_in62,local6_out62,
local6_in63,local6_out63,
local6_in64,local6_out64,
local6_in65,local6_out65,
local6_in66,local6_out66,
local6_in67,local6_out67,
local6_in68,local6_out68,
local6_in69,local6_out69,
local7_in70,local7_out70,
local7_in71,local7_out71,
local7_in72,local7_out72,
local7_in73,local7_out73,
local7_in74,local7_out74,
local7_in75,local7_out75,
local7_in76,local7_out76,
local7_in77,local7_out77,
local7_in78,local7_out78,
local7_in79,local7_out79,
local8_in80,local8_out80,
local8_in81,local8_out81,
local8_in82,local8_out82,
local8_in83,local8_out83,
local8_in84,local8_out84,
local8_in85,local8_out85,
local8_in86,local8_out86,
local8_in87,local8_out87,
local8_in88,local8_out88,
local8_in89,local8_out89,
local9_in90,local9_out90,
local9_in91,local9_out91,
local9_in92,local9_out92,
local9_in93,local9_out93,
local9_in94,local9_out94,
local9_in95,local9_out95,
local9_in96,local9_out96,
local9_in97,local9_out97,
local9_in98,local9_out98,
local9_in99,local9_out99,
clk, reset,  Write, Read);
input clk, reset, Write, Read; 
parameter DATAWID = 32;
input [DATAWID-1:0] local0_in00;
output [DATAWID-1:0] local0_out00;
input [DATAWID-1:0] local0_in01;
output [DATAWID-1:0] local0_out01;
input [DATAWID-1:0] local0_in02;
output [DATAWID-1:0] local0_out02;
input [DATAWID-1:0] local0_in03;
output [DATAWID-1:0] local0_out03;
input [DATAWID-1:0] local0_in04;
output [DATAWID-1:0] local0_out04;
input [DATAWID-1:0] local0_in05;
output [DATAWID-1:0] local0_out05;
input [DATAWID-1:0] local0_in06;
output [DATAWID-1:0] local0_out06;
input [DATAWID-1:0] local0_in07;
output [DATAWID-1:0] local0_out07;
input [DATAWID-1:0] local0_in08;
output [DATAWID-1:0] local0_out08;
input [DATAWID-1:0] local0_in09;
output [DATAWID-1:0] local0_out09;
input [DATAWID-1:0] local1_in10;
output [DATAWID-1:0] local1_out10;
input [DATAWID-1:0] local1_in11;
output [DATAWID-1:0] local1_out11;
input [DATAWID-1:0] local1_in12;
output [DATAWID-1:0] local1_out12;
input [DATAWID-1:0] local1_in13;
output [DATAWID-1:0] local1_out13;
input [DATAWID-1:0] local1_in14;
output [DATAWID-1:0] local1_out14;
input [DATAWID-1:0] local1_in15;
output [DATAWID-1:0] local1_out15;
input [DATAWID-1:0] local1_in16;
output [DATAWID-1:0] local1_out16;
input [DATAWID-1:0] local1_in17;
output [DATAWID-1:0] local1_out17;
input [DATAWID-1:0] local1_in18;
output [DATAWID-1:0] local1_out18;
input [DATAWID-1:0] local1_in19;
output [DATAWID-1:0] local1_out19;
input [DATAWID-1:0] local2_in20;
output [DATAWID-1:0] local2_out20;
input [DATAWID-1:0] local2_in21;
output [DATAWID-1:0] local2_out21;
input [DATAWID-1:0] local2_in22;
output [DATAWID-1:0] local2_out22;
input [DATAWID-1:0] local2_in23;
output [DATAWID-1:0] local2_out23;
input [DATAWID-1:0] local2_in24;
output [DATAWID-1:0] local2_out24;
input [DATAWID-1:0] local2_in25;
output [DATAWID-1:0] local2_out25;
input [DATAWID-1:0] local2_in26;
output [DATAWID-1:0] local2_out26;
input [DATAWID-1:0] local2_in27;
output [DATAWID-1:0] local2_out27;
input [DATAWID-1:0] local2_in28;
output [DATAWID-1:0] local2_out28;
input [DATAWID-1:0] local2_in29;
output [DATAWID-1:0] local2_out29;
input [DATAWID-1:0] local3_in30;
output [DATAWID-1:0] local3_out30;
input [DATAWID-1:0] local3_in31;
output [DATAWID-1:0] local3_out31;
input [DATAWID-1:0] local3_in32;
output [DATAWID-1:0] local3_out32;
input [DATAWID-1:0] local3_in33;
output [DATAWID-1:0] local3_out33;
input [DATAWID-1:0] local3_in34;
output [DATAWID-1:0] local3_out34;
input [DATAWID-1:0] local3_in35;
output [DATAWID-1:0] local3_out35;
input [DATAWID-1:0] local3_in36;
output [DATAWID-1:0] local3_out36;
input [DATAWID-1:0] local3_in37;
output [DATAWID-1:0] local3_out37;
input [DATAWID-1:0] local3_in38;
output [DATAWID-1:0] local3_out38;
input [DATAWID-1:0] local3_in39;
output [DATAWID-1:0] local3_out39;
input [DATAWID-1:0] local4_in40;
output [DATAWID-1:0] local4_out40;
input [DATAWID-1:0] local4_in41;
output [DATAWID-1:0] local4_out41;
input [DATAWID-1:0] local4_in42;
output [DATAWID-1:0] local4_out42;
input [DATAWID-1:0] local4_in43;
output [DATAWID-1:0] local4_out43;
input [DATAWID-1:0] local4_in44;
output [DATAWID-1:0] local4_out44;
input [DATAWID-1:0] local4_in45;
output [DATAWID-1:0] local4_out45;
input [DATAWID-1:0] local4_in46;
output [DATAWID-1:0] local4_out46;
input [DATAWID-1:0] local4_in47;
output [DATAWID-1:0] local4_out47;
input [DATAWID-1:0] local4_in48;
output [DATAWID-1:0] local4_out48;
input [DATAWID-1:0] local4_in49;
output [DATAWID-1:0] local4_out49;
input [DATAWID-1:0] local5_in50;
output [DATAWID-1:0] local5_out50;
input [DATAWID-1:0] local5_in51;
output [DATAWID-1:0] local5_out51;
input [DATAWID-1:0] local5_in52;
output [DATAWID-1:0] local5_out52;
input [DATAWID-1:0] local5_in53;
output [DATAWID-1:0] local5_out53;
input [DATAWID-1:0] local5_in54;
output [DATAWID-1:0] local5_out54;
input [DATAWID-1:0] local5_in55;
output [DATAWID-1:0] local5_out55;
input [DATAWID-1:0] local5_in56;
output [DATAWID-1:0] local5_out56;
input [DATAWID-1:0] local5_in57;
output [DATAWID-1:0] local5_out57;
input [DATAWID-1:0] local5_in58;
output [DATAWID-1:0] local5_out58;
input [DATAWID-1:0] local5_in59;
output [DATAWID-1:0] local5_out59;
input [DATAWID-1:0] local6_in60;
output [DATAWID-1:0] local6_out60;
input [DATAWID-1:0] local6_in61;
output [DATAWID-1:0] local6_out61;
input [DATAWID-1:0] local6_in62;
output [DATAWID-1:0] local6_out62;
input [DATAWID-1:0] local6_in63;
output [DATAWID-1:0] local6_out63;
input [DATAWID-1:0] local6_in64;
output [DATAWID-1:0] local6_out64;
input [DATAWID-1:0] local6_in65;
output [DATAWID-1:0] local6_out65;
input [DATAWID-1:0] local6_in66;
output [DATAWID-1:0] local6_out66;
input [DATAWID-1:0] local6_in67;
output [DATAWID-1:0] local6_out67;
input [DATAWID-1:0] local6_in68;
output [DATAWID-1:0] local6_out68;
input [DATAWID-1:0] local6_in69;
output [DATAWID-1:0] local6_out69;
input [DATAWID-1:0] local7_in70;
output [DATAWID-1:0] local7_out70;
input [DATAWID-1:0] local7_in71;
output [DATAWID-1:0] local7_out71;
input [DATAWID-1:0] local7_in72;
output [DATAWID-1:0] local7_out72;
input [DATAWID-1:0] local7_in73;
output [DATAWID-1:0] local7_out73;
input [DATAWID-1:0] local7_in74;
output [DATAWID-1:0] local7_out74;
input [DATAWID-1:0] local7_in75;
output [DATAWID-1:0] local7_out75;
input [DATAWID-1:0] local7_in76;
output [DATAWID-1:0] local7_out76;
input [DATAWID-1:0] local7_in77;
output [DATAWID-1:0] local7_out77;
input [DATAWID-1:0] local7_in78;
output [DATAWID-1:0] local7_out78;
input [DATAWID-1:0] local7_in79;
output [DATAWID-1:0] local7_out79;
input [DATAWID-1:0] local8_in80;
output [DATAWID-1:0] local8_out80;
input [DATAWID-1:0] local8_in81;
output [DATAWID-1:0] local8_out81;
input [DATAWID-1:0] local8_in82;
output [DATAWID-1:0] local8_out82;
input [DATAWID-1:0] local8_in83;
output [DATAWID-1:0] local8_out83;
input [DATAWID-1:0] local8_in84;
output [DATAWID-1:0] local8_out84;
input [DATAWID-1:0] local8_in85;
output [DATAWID-1:0] local8_out85;
input [DATAWID-1:0] local8_in86;
output [DATAWID-1:0] local8_out86;
input [DATAWID-1:0] local8_in87;
output [DATAWID-1:0] local8_out87;
input [DATAWID-1:0] local8_in88;
output [DATAWID-1:0] local8_out88;
input [DATAWID-1:0] local8_in89;
output [DATAWID-1:0] local8_out89;
input [DATAWID-1:0] local9_in90;
output [DATAWID-1:0] local9_out90;
input [DATAWID-1:0] local9_in91;
output [DATAWID-1:0] local9_out91;
input [DATAWID-1:0] local9_in92;
output [DATAWID-1:0] local9_out92;
input [DATAWID-1:0] local9_in93;
output [DATAWID-1:0] local9_out93;
input [DATAWID-1:0] local9_in94;
output [DATAWID-1:0] local9_out94;
input [DATAWID-1:0] local9_in95;
output [DATAWID-1:0] local9_out95;
input [DATAWID-1:0] local9_in96;
output [DATAWID-1:0] local9_out96;
input [DATAWID-1:0] local9_in97;
output [DATAWID-1:0] local9_out97;
input [DATAWID-1:0] local9_in98;
output [DATAWID-1:0] local9_out98;
input [DATAWID-1:0] local9_in99;
output [DATAWID-1:0] local9_out99;
reg [DATAWID-1:0] east0_in00;
reg [DATAWID-1:0] west0_in00;
reg [DATAWID-1:0] north0_in00;
reg [DATAWID-1:0] south0_in00;
reg [DATAWID-1:0] east0_in01;
reg [DATAWID-1:0] west0_in01;
reg [DATAWID-1:0] north0_in01;
reg [DATAWID-1:0] south0_in01;
reg [DATAWID-1:0] east0_in02;
reg [DATAWID-1:0] west0_in02;
reg [DATAWID-1:0] north0_in02;
reg [DATAWID-1:0] south0_in02;
reg [DATAWID-1:0] east0_in03;
reg [DATAWID-1:0] west0_in03;
reg [DATAWID-1:0] north0_in03;
reg [DATAWID-1:0] south0_in03;
reg [DATAWID-1:0] east0_in04;
reg [DATAWID-1:0] west0_in04;
reg [DATAWID-1:0] north0_in04;
reg [DATAWID-1:0] south0_in04;
reg [DATAWID-1:0] east0_in05;
reg [DATAWID-1:0] west0_in05;
reg [DATAWID-1:0] north0_in05;
reg [DATAWID-1:0] south0_in05;
reg [DATAWID-1:0] east0_in06;
reg [DATAWID-1:0] west0_in06;
reg [DATAWID-1:0] north0_in06;
reg [DATAWID-1:0] south0_in06;
reg [DATAWID-1:0] east0_in07;
reg [DATAWID-1:0] west0_in07;
reg [DATAWID-1:0] north0_in07;
reg [DATAWID-1:0] south0_in07;
reg [DATAWID-1:0] east0_in08;
reg [DATAWID-1:0] west0_in08;
reg [DATAWID-1:0] north0_in08;
reg [DATAWID-1:0] south0_in08;
reg [DATAWID-1:0] east0_in09;
reg [DATAWID-1:0] west0_in09;
reg [DATAWID-1:0] north0_in09;
reg [DATAWID-1:0] south0_in09;
reg [DATAWID-1:0] east1_in10;
reg [DATAWID-1:0] west1_in10;
reg [DATAWID-1:0] north1_in10;
reg [DATAWID-1:0] south1_in10;
reg [DATAWID-1:0] east1_in11;
reg [DATAWID-1:0] west1_in11;
reg [DATAWID-1:0] north1_in11;
reg [DATAWID-1:0] south1_in11;
reg [DATAWID-1:0] east1_in12;
reg [DATAWID-1:0] west1_in12;
reg [DATAWID-1:0] north1_in12;
reg [DATAWID-1:0] south1_in12;
reg [DATAWID-1:0] east1_in13;
reg [DATAWID-1:0] west1_in13;
reg [DATAWID-1:0] north1_in13;
reg [DATAWID-1:0] south1_in13;
reg [DATAWID-1:0] east1_in14;
reg [DATAWID-1:0] west1_in14;
reg [DATAWID-1:0] north1_in14;
reg [DATAWID-1:0] south1_in14;
reg [DATAWID-1:0] east1_in15;
reg [DATAWID-1:0] west1_in15;
reg [DATAWID-1:0] north1_in15;
reg [DATAWID-1:0] south1_in15;
reg [DATAWID-1:0] east1_in16;
reg [DATAWID-1:0] west1_in16;
reg [DATAWID-1:0] north1_in16;
reg [DATAWID-1:0] south1_in16;
reg [DATAWID-1:0] east1_in17;
reg [DATAWID-1:0] west1_in17;
reg [DATAWID-1:0] north1_in17;
reg [DATAWID-1:0] south1_in17;
reg [DATAWID-1:0] east1_in18;
reg [DATAWID-1:0] west1_in18;
reg [DATAWID-1:0] north1_in18;
reg [DATAWID-1:0] south1_in18;
reg [DATAWID-1:0] east1_in19;
reg [DATAWID-1:0] west1_in19;
reg [DATAWID-1:0] north1_in19;
reg [DATAWID-1:0] south1_in19;
reg [DATAWID-1:0] east2_in20;
reg [DATAWID-1:0] west2_in20;
reg [DATAWID-1:0] north2_in20;
reg [DATAWID-1:0] south2_in20;
reg [DATAWID-1:0] east2_in21;
reg [DATAWID-1:0] west2_in21;
reg [DATAWID-1:0] north2_in21;
reg [DATAWID-1:0] south2_in21;
reg [DATAWID-1:0] east2_in22;
reg [DATAWID-1:0] west2_in22;
reg [DATAWID-1:0] north2_in22;
reg [DATAWID-1:0] south2_in22;
reg [DATAWID-1:0] east2_in23;
reg [DATAWID-1:0] west2_in23;
reg [DATAWID-1:0] north2_in23;
reg [DATAWID-1:0] south2_in23;
reg [DATAWID-1:0] east2_in24;
reg [DATAWID-1:0] west2_in24;
reg [DATAWID-1:0] north2_in24;
reg [DATAWID-1:0] south2_in24;
reg [DATAWID-1:0] east2_in25;
reg [DATAWID-1:0] west2_in25;
reg [DATAWID-1:0] north2_in25;
reg [DATAWID-1:0] south2_in25;
reg [DATAWID-1:0] east2_in26;
reg [DATAWID-1:0] west2_in26;
reg [DATAWID-1:0] north2_in26;
reg [DATAWID-1:0] south2_in26;
reg [DATAWID-1:0] east2_in27;
reg [DATAWID-1:0] west2_in27;
reg [DATAWID-1:0] north2_in27;
reg [DATAWID-1:0] south2_in27;
reg [DATAWID-1:0] east2_in28;
reg [DATAWID-1:0] west2_in28;
reg [DATAWID-1:0] north2_in28;
reg [DATAWID-1:0] south2_in28;
reg [DATAWID-1:0] east2_in29;
reg [DATAWID-1:0] west2_in29;
reg [DATAWID-1:0] north2_in29;
reg [DATAWID-1:0] south2_in29;
reg [DATAWID-1:0] east3_in30;
reg [DATAWID-1:0] west3_in30;
reg [DATAWID-1:0] north3_in30;
reg [DATAWID-1:0] south3_in30;
reg [DATAWID-1:0] east3_in31;
reg [DATAWID-1:0] west3_in31;
reg [DATAWID-1:0] north3_in31;
reg [DATAWID-1:0] south3_in31;
reg [DATAWID-1:0] east3_in32;
reg [DATAWID-1:0] west3_in32;
reg [DATAWID-1:0] north3_in32;
reg [DATAWID-1:0] south3_in32;
reg [DATAWID-1:0] east3_in33;
reg [DATAWID-1:0] west3_in33;
reg [DATAWID-1:0] north3_in33;
reg [DATAWID-1:0] south3_in33;
reg [DATAWID-1:0] east3_in34;
reg [DATAWID-1:0] west3_in34;
reg [DATAWID-1:0] north3_in34;
reg [DATAWID-1:0] south3_in34;
reg [DATAWID-1:0] east3_in35;
reg [DATAWID-1:0] west3_in35;
reg [DATAWID-1:0] north3_in35;
reg [DATAWID-1:0] south3_in35;
reg [DATAWID-1:0] east3_in36;
reg [DATAWID-1:0] west3_in36;
reg [DATAWID-1:0] north3_in36;
reg [DATAWID-1:0] south3_in36;
reg [DATAWID-1:0] east3_in37;
reg [DATAWID-1:0] west3_in37;
reg [DATAWID-1:0] north3_in37;
reg [DATAWID-1:0] south3_in37;
reg [DATAWID-1:0] east3_in38;
reg [DATAWID-1:0] west3_in38;
reg [DATAWID-1:0] north3_in38;
reg [DATAWID-1:0] south3_in38;
reg [DATAWID-1:0] east3_in39;
reg [DATAWID-1:0] west3_in39;
reg [DATAWID-1:0] north3_in39;
reg [DATAWID-1:0] south3_in39;
reg [DATAWID-1:0] east4_in40;
reg [DATAWID-1:0] west4_in40;
reg [DATAWID-1:0] north4_in40;
reg [DATAWID-1:0] south4_in40;
reg [DATAWID-1:0] east4_in41;
reg [DATAWID-1:0] west4_in41;
reg [DATAWID-1:0] north4_in41;
reg [DATAWID-1:0] south4_in41;
reg [DATAWID-1:0] east4_in42;
reg [DATAWID-1:0] west4_in42;
reg [DATAWID-1:0] north4_in42;
reg [DATAWID-1:0] south4_in42;
reg [DATAWID-1:0] east4_in43;
reg [DATAWID-1:0] west4_in43;
reg [DATAWID-1:0] north4_in43;
reg [DATAWID-1:0] south4_in43;
reg [DATAWID-1:0] east4_in44;
reg [DATAWID-1:0] west4_in44;
reg [DATAWID-1:0] north4_in44;
reg [DATAWID-1:0] south4_in44;
reg [DATAWID-1:0] east4_in45;
reg [DATAWID-1:0] west4_in45;
reg [DATAWID-1:0] north4_in45;
reg [DATAWID-1:0] south4_in45;
reg [DATAWID-1:0] east4_in46;
reg [DATAWID-1:0] west4_in46;
reg [DATAWID-1:0] north4_in46;
reg [DATAWID-1:0] south4_in46;
reg [DATAWID-1:0] east4_in47;
reg [DATAWID-1:0] west4_in47;
reg [DATAWID-1:0] north4_in47;
reg [DATAWID-1:0] south4_in47;
reg [DATAWID-1:0] east4_in48;
reg [DATAWID-1:0] west4_in48;
reg [DATAWID-1:0] north4_in48;
reg [DATAWID-1:0] south4_in48;
reg [DATAWID-1:0] east4_in49;
reg [DATAWID-1:0] west4_in49;
reg [DATAWID-1:0] north4_in49;
reg [DATAWID-1:0] south4_in49;
reg [DATAWID-1:0] east5_in50;
reg [DATAWID-1:0] west5_in50;
reg [DATAWID-1:0] north5_in50;
reg [DATAWID-1:0] south5_in50;
reg [DATAWID-1:0] east5_in51;
reg [DATAWID-1:0] west5_in51;
reg [DATAWID-1:0] north5_in51;
reg [DATAWID-1:0] south5_in51;
reg [DATAWID-1:0] east5_in52;
reg [DATAWID-1:0] west5_in52;
reg [DATAWID-1:0] north5_in52;
reg [DATAWID-1:0] south5_in52;
reg [DATAWID-1:0] east5_in53;
reg [DATAWID-1:0] west5_in53;
reg [DATAWID-1:0] north5_in53;
reg [DATAWID-1:0] south5_in53;
reg [DATAWID-1:0] east5_in54;
reg [DATAWID-1:0] west5_in54;
reg [DATAWID-1:0] north5_in54;
reg [DATAWID-1:0] south5_in54;
reg [DATAWID-1:0] east5_in55;
reg [DATAWID-1:0] west5_in55;
reg [DATAWID-1:0] north5_in55;
reg [DATAWID-1:0] south5_in55;
reg [DATAWID-1:0] east5_in56;
reg [DATAWID-1:0] west5_in56;
reg [DATAWID-1:0] north5_in56;
reg [DATAWID-1:0] south5_in56;
reg [DATAWID-1:0] east5_in57;
reg [DATAWID-1:0] west5_in57;
reg [DATAWID-1:0] north5_in57;
reg [DATAWID-1:0] south5_in57;
reg [DATAWID-1:0] east5_in58;
reg [DATAWID-1:0] west5_in58;
reg [DATAWID-1:0] north5_in58;
reg [DATAWID-1:0] south5_in58;
reg [DATAWID-1:0] east5_in59;
reg [DATAWID-1:0] west5_in59;
reg [DATAWID-1:0] north5_in59;
reg [DATAWID-1:0] south5_in59;
reg [DATAWID-1:0] east6_in60;
reg [DATAWID-1:0] west6_in60;
reg [DATAWID-1:0] north6_in60;
reg [DATAWID-1:0] south6_in60;
reg [DATAWID-1:0] east6_in61;
reg [DATAWID-1:0] west6_in61;
reg [DATAWID-1:0] north6_in61;
reg [DATAWID-1:0] south6_in61;
reg [DATAWID-1:0] east6_in62;
reg [DATAWID-1:0] west6_in62;
reg [DATAWID-1:0] north6_in62;
reg [DATAWID-1:0] south6_in62;
reg [DATAWID-1:0] east6_in63;
reg [DATAWID-1:0] west6_in63;
reg [DATAWID-1:0] north6_in63;
reg [DATAWID-1:0] south6_in63;
reg [DATAWID-1:0] east6_in64;
reg [DATAWID-1:0] west6_in64;
reg [DATAWID-1:0] north6_in64;
reg [DATAWID-1:0] south6_in64;
reg [DATAWID-1:0] east6_in65;
reg [DATAWID-1:0] west6_in65;
reg [DATAWID-1:0] north6_in65;
reg [DATAWID-1:0] south6_in65;
reg [DATAWID-1:0] east6_in66;
reg [DATAWID-1:0] west6_in66;
reg [DATAWID-1:0] north6_in66;
reg [DATAWID-1:0] south6_in66;
reg [DATAWID-1:0] east6_in67;
reg [DATAWID-1:0] west6_in67;
reg [DATAWID-1:0] north6_in67;
reg [DATAWID-1:0] south6_in67;
reg [DATAWID-1:0] east6_in68;
reg [DATAWID-1:0] west6_in68;
reg [DATAWID-1:0] north6_in68;
reg [DATAWID-1:0] south6_in68;
reg [DATAWID-1:0] east6_in69;
reg [DATAWID-1:0] west6_in69;
reg [DATAWID-1:0] north6_in69;
reg [DATAWID-1:0] south6_in69;
reg [DATAWID-1:0] east7_in70;
reg [DATAWID-1:0] west7_in70;
reg [DATAWID-1:0] north7_in70;
reg [DATAWID-1:0] south7_in70;
reg [DATAWID-1:0] east7_in71;
reg [DATAWID-1:0] west7_in71;
reg [DATAWID-1:0] north7_in71;
reg [DATAWID-1:0] south7_in71;
reg [DATAWID-1:0] east7_in72;
reg [DATAWID-1:0] west7_in72;
reg [DATAWID-1:0] north7_in72;
reg [DATAWID-1:0] south7_in72;
reg [DATAWID-1:0] east7_in73;
reg [DATAWID-1:0] west7_in73;
reg [DATAWID-1:0] north7_in73;
reg [DATAWID-1:0] south7_in73;
reg [DATAWID-1:0] east7_in74;
reg [DATAWID-1:0] west7_in74;
reg [DATAWID-1:0] north7_in74;
reg [DATAWID-1:0] south7_in74;
reg [DATAWID-1:0] east7_in75;
reg [DATAWID-1:0] west7_in75;
reg [DATAWID-1:0] north7_in75;
reg [DATAWID-1:0] south7_in75;
reg [DATAWID-1:0] east7_in76;
reg [DATAWID-1:0] west7_in76;
reg [DATAWID-1:0] north7_in76;
reg [DATAWID-1:0] south7_in76;
reg [DATAWID-1:0] east7_in77;
reg [DATAWID-1:0] west7_in77;
reg [DATAWID-1:0] north7_in77;
reg [DATAWID-1:0] south7_in77;
reg [DATAWID-1:0] east7_in78;
reg [DATAWID-1:0] west7_in78;
reg [DATAWID-1:0] north7_in78;
reg [DATAWID-1:0] south7_in78;
reg [DATAWID-1:0] east7_in79;
reg [DATAWID-1:0] west7_in79;
reg [DATAWID-1:0] north7_in79;
reg [DATAWID-1:0] south7_in79;
reg [DATAWID-1:0] east8_in80;
reg [DATAWID-1:0] west8_in80;
reg [DATAWID-1:0] north8_in80;
reg [DATAWID-1:0] south8_in80;
reg [DATAWID-1:0] east8_in81;
reg [DATAWID-1:0] west8_in81;
reg [DATAWID-1:0] north8_in81;
reg [DATAWID-1:0] south8_in81;
reg [DATAWID-1:0] east8_in82;
reg [DATAWID-1:0] west8_in82;
reg [DATAWID-1:0] north8_in82;
reg [DATAWID-1:0] south8_in82;
reg [DATAWID-1:0] east8_in83;
reg [DATAWID-1:0] west8_in83;
reg [DATAWID-1:0] north8_in83;
reg [DATAWID-1:0] south8_in83;
reg [DATAWID-1:0] east8_in84;
reg [DATAWID-1:0] west8_in84;
reg [DATAWID-1:0] north8_in84;
reg [DATAWID-1:0] south8_in84;
reg [DATAWID-1:0] east8_in85;
reg [DATAWID-1:0] west8_in85;
reg [DATAWID-1:0] north8_in85;
reg [DATAWID-1:0] south8_in85;
reg [DATAWID-1:0] east8_in86;
reg [DATAWID-1:0] west8_in86;
reg [DATAWID-1:0] north8_in86;
reg [DATAWID-1:0] south8_in86;
reg [DATAWID-1:0] east8_in87;
reg [DATAWID-1:0] west8_in87;
reg [DATAWID-1:0] north8_in87;
reg [DATAWID-1:0] south8_in87;
reg [DATAWID-1:0] east8_in88;
reg [DATAWID-1:0] west8_in88;
reg [DATAWID-1:0] north8_in88;
reg [DATAWID-1:0] south8_in88;
reg [DATAWID-1:0] east8_in89;
reg [DATAWID-1:0] west8_in89;
reg [DATAWID-1:0] north8_in89;
reg [DATAWID-1:0] south8_in89;
reg [DATAWID-1:0] east9_in90;
reg [DATAWID-1:0] west9_in90;
reg [DATAWID-1:0] north9_in90;
reg [DATAWID-1:0] south9_in90;
reg [DATAWID-1:0] east9_in91;
reg [DATAWID-1:0] west9_in91;
reg [DATAWID-1:0] north9_in91;
reg [DATAWID-1:0] south9_in91;
reg [DATAWID-1:0] east9_in92;
reg [DATAWID-1:0] west9_in92;
reg [DATAWID-1:0] north9_in92;
reg [DATAWID-1:0] south9_in92;
reg [DATAWID-1:0] east9_in93;
reg [DATAWID-1:0] west9_in93;
reg [DATAWID-1:0] north9_in93;
reg [DATAWID-1:0] south9_in93;
reg [DATAWID-1:0] east9_in94;
reg [DATAWID-1:0] west9_in94;
reg [DATAWID-1:0] north9_in94;
reg [DATAWID-1:0] south9_in94;
reg [DATAWID-1:0] east9_in95;
reg [DATAWID-1:0] west9_in95;
reg [DATAWID-1:0] north9_in95;
reg [DATAWID-1:0] south9_in95;
reg [DATAWID-1:0] east9_in96;
reg [DATAWID-1:0] west9_in96;
reg [DATAWID-1:0] north9_in96;
reg [DATAWID-1:0] south9_in96;
reg [DATAWID-1:0] east9_in97;
reg [DATAWID-1:0] west9_in97;
reg [DATAWID-1:0] north9_in97;
reg [DATAWID-1:0] south9_in97;
reg [DATAWID-1:0] east9_in98;
reg [DATAWID-1:0] west9_in98;
reg [DATAWID-1:0] north9_in98;
reg [DATAWID-1:0] south9_in98;
reg [DATAWID-1:0] east9_in99;
reg [DATAWID-1:0] west9_in99;
reg [DATAWID-1:0] north9_in99;
reg [DATAWID-1:0] south9_in99;
wire [DATAWID-1:0] east0_out00;
wire [DATAWID-1:0] west0_out00;
wire [DATAWID-1:0] north0_out00;
wire [DATAWID-1:0] south0_out00;
wire [DATAWID-1:0] east0_out01;
wire [DATAWID-1:0] west0_out01;
wire [DATAWID-1:0] north0_out01;
wire [DATAWID-1:0] south0_out01;
wire [DATAWID-1:0] east0_out02;
wire [DATAWID-1:0] west0_out02;
wire [DATAWID-1:0] north0_out02;
wire [DATAWID-1:0] south0_out02;
wire [DATAWID-1:0] east0_out03;
wire [DATAWID-1:0] west0_out03;
wire [DATAWID-1:0] north0_out03;
wire [DATAWID-1:0] south0_out03;
wire [DATAWID-1:0] east0_out04;
wire [DATAWID-1:0] west0_out04;
wire [DATAWID-1:0] north0_out04;
wire [DATAWID-1:0] south0_out04;
wire [DATAWID-1:0] east0_out05;
wire [DATAWID-1:0] west0_out05;
wire [DATAWID-1:0] north0_out05;
wire [DATAWID-1:0] south0_out05;
wire [DATAWID-1:0] east0_out06;
wire [DATAWID-1:0] west0_out06;
wire [DATAWID-1:0] north0_out06;
wire [DATAWID-1:0] south0_out06;
wire [DATAWID-1:0] east0_out07;
wire [DATAWID-1:0] west0_out07;
wire [DATAWID-1:0] north0_out07;
wire [DATAWID-1:0] south0_out07;
wire [DATAWID-1:0] east0_out08;
wire [DATAWID-1:0] west0_out08;
wire [DATAWID-1:0] north0_out08;
wire [DATAWID-1:0] south0_out08;
wire [DATAWID-1:0] east0_out09;
wire [DATAWID-1:0] west0_out09;
wire [DATAWID-1:0] north0_out09;
wire [DATAWID-1:0] south0_out09;
wire [DATAWID-1:0] east1_out10;
wire [DATAWID-1:0] west1_out10;
wire [DATAWID-1:0] north1_out10;
wire [DATAWID-1:0] south1_out10;
wire [DATAWID-1:0] east1_out11;
wire [DATAWID-1:0] west1_out11;
wire [DATAWID-1:0] north1_out11;
wire [DATAWID-1:0] south1_out11;
wire [DATAWID-1:0] east1_out12;
wire [DATAWID-1:0] west1_out12;
wire [DATAWID-1:0] north1_out12;
wire [DATAWID-1:0] south1_out12;
wire [DATAWID-1:0] east1_out13;
wire [DATAWID-1:0] west1_out13;
wire [DATAWID-1:0] north1_out13;
wire [DATAWID-1:0] south1_out13;
wire [DATAWID-1:0] east1_out14;
wire [DATAWID-1:0] west1_out14;
wire [DATAWID-1:0] north1_out14;
wire [DATAWID-1:0] south1_out14;
wire [DATAWID-1:0] east1_out15;
wire [DATAWID-1:0] west1_out15;
wire [DATAWID-1:0] north1_out15;
wire [DATAWID-1:0] south1_out15;
wire [DATAWID-1:0] east1_out16;
wire [DATAWID-1:0] west1_out16;
wire [DATAWID-1:0] north1_out16;
wire [DATAWID-1:0] south1_out16;
wire [DATAWID-1:0] east1_out17;
wire [DATAWID-1:0] west1_out17;
wire [DATAWID-1:0] north1_out17;
wire [DATAWID-1:0] south1_out17;
wire [DATAWID-1:0] east1_out18;
wire [DATAWID-1:0] west1_out18;
wire [DATAWID-1:0] north1_out18;
wire [DATAWID-1:0] south1_out18;
wire [DATAWID-1:0] east1_out19;
wire [DATAWID-1:0] west1_out19;
wire [DATAWID-1:0] north1_out19;
wire [DATAWID-1:0] south1_out19;
wire [DATAWID-1:0] east2_out20;
wire [DATAWID-1:0] west2_out20;
wire [DATAWID-1:0] north2_out20;
wire [DATAWID-1:0] south2_out20;
wire [DATAWID-1:0] east2_out21;
wire [DATAWID-1:0] west2_out21;
wire [DATAWID-1:0] north2_out21;
wire [DATAWID-1:0] south2_out21;
wire [DATAWID-1:0] east2_out22;
wire [DATAWID-1:0] west2_out22;
wire [DATAWID-1:0] north2_out22;
wire [DATAWID-1:0] south2_out22;
wire [DATAWID-1:0] east2_out23;
wire [DATAWID-1:0] west2_out23;
wire [DATAWID-1:0] north2_out23;
wire [DATAWID-1:0] south2_out23;
wire [DATAWID-1:0] east2_out24;
wire [DATAWID-1:0] west2_out24;
wire [DATAWID-1:0] north2_out24;
wire [DATAWID-1:0] south2_out24;
wire [DATAWID-1:0] east2_out25;
wire [DATAWID-1:0] west2_out25;
wire [DATAWID-1:0] north2_out25;
wire [DATAWID-1:0] south2_out25;
wire [DATAWID-1:0] east2_out26;
wire [DATAWID-1:0] west2_out26;
wire [DATAWID-1:0] north2_out26;
wire [DATAWID-1:0] south2_out26;
wire [DATAWID-1:0] east2_out27;
wire [DATAWID-1:0] west2_out27;
wire [DATAWID-1:0] north2_out27;
wire [DATAWID-1:0] south2_out27;
wire [DATAWID-1:0] east2_out28;
wire [DATAWID-1:0] west2_out28;
wire [DATAWID-1:0] north2_out28;
wire [DATAWID-1:0] south2_out28;
wire [DATAWID-1:0] east2_out29;
wire [DATAWID-1:0] west2_out29;
wire [DATAWID-1:0] north2_out29;
wire [DATAWID-1:0] south2_out29;
wire [DATAWID-1:0] east3_out30;
wire [DATAWID-1:0] west3_out30;
wire [DATAWID-1:0] north3_out30;
wire [DATAWID-1:0] south3_out30;
wire [DATAWID-1:0] east3_out31;
wire [DATAWID-1:0] west3_out31;
wire [DATAWID-1:0] north3_out31;
wire [DATAWID-1:0] south3_out31;
wire [DATAWID-1:0] east3_out32;
wire [DATAWID-1:0] west3_out32;
wire [DATAWID-1:0] north3_out32;
wire [DATAWID-1:0] south3_out32;
wire [DATAWID-1:0] east3_out33;
wire [DATAWID-1:0] west3_out33;
wire [DATAWID-1:0] north3_out33;
wire [DATAWID-1:0] south3_out33;
wire [DATAWID-1:0] east3_out34;
wire [DATAWID-1:0] west3_out34;
wire [DATAWID-1:0] north3_out34;
wire [DATAWID-1:0] south3_out34;
wire [DATAWID-1:0] east3_out35;
wire [DATAWID-1:0] west3_out35;
wire [DATAWID-1:0] north3_out35;
wire [DATAWID-1:0] south3_out35;
wire [DATAWID-1:0] east3_out36;
wire [DATAWID-1:0] west3_out36;
wire [DATAWID-1:0] north3_out36;
wire [DATAWID-1:0] south3_out36;
wire [DATAWID-1:0] east3_out37;
wire [DATAWID-1:0] west3_out37;
wire [DATAWID-1:0] north3_out37;
wire [DATAWID-1:0] south3_out37;
wire [DATAWID-1:0] east3_out38;
wire [DATAWID-1:0] west3_out38;
wire [DATAWID-1:0] north3_out38;
wire [DATAWID-1:0] south3_out38;
wire [DATAWID-1:0] east3_out39;
wire [DATAWID-1:0] west3_out39;
wire [DATAWID-1:0] north3_out39;
wire [DATAWID-1:0] south3_out39;
wire [DATAWID-1:0] east4_out40;
wire [DATAWID-1:0] west4_out40;
wire [DATAWID-1:0] north4_out40;
wire [DATAWID-1:0] south4_out40;
wire [DATAWID-1:0] east4_out41;
wire [DATAWID-1:0] west4_out41;
wire [DATAWID-1:0] north4_out41;
wire [DATAWID-1:0] south4_out41;
wire [DATAWID-1:0] east4_out42;
wire [DATAWID-1:0] west4_out42;
wire [DATAWID-1:0] north4_out42;
wire [DATAWID-1:0] south4_out42;
wire [DATAWID-1:0] east4_out43;
wire [DATAWID-1:0] west4_out43;
wire [DATAWID-1:0] north4_out43;
wire [DATAWID-1:0] south4_out43;
wire [DATAWID-1:0] east4_out44;
wire [DATAWID-1:0] west4_out44;
wire [DATAWID-1:0] north4_out44;
wire [DATAWID-1:0] south4_out44;
wire [DATAWID-1:0] east4_out45;
wire [DATAWID-1:0] west4_out45;
wire [DATAWID-1:0] north4_out45;
wire [DATAWID-1:0] south4_out45;
wire [DATAWID-1:0] east4_out46;
wire [DATAWID-1:0] west4_out46;
wire [DATAWID-1:0] north4_out46;
wire [DATAWID-1:0] south4_out46;
wire [DATAWID-1:0] east4_out47;
wire [DATAWID-1:0] west4_out47;
wire [DATAWID-1:0] north4_out47;
wire [DATAWID-1:0] south4_out47;
wire [DATAWID-1:0] east4_out48;
wire [DATAWID-1:0] west4_out48;
wire [DATAWID-1:0] north4_out48;
wire [DATAWID-1:0] south4_out48;
wire [DATAWID-1:0] east4_out49;
wire [DATAWID-1:0] west4_out49;
wire [DATAWID-1:0] north4_out49;
wire [DATAWID-1:0] south4_out49;
wire [DATAWID-1:0] east5_out50;
wire [DATAWID-1:0] west5_out50;
wire [DATAWID-1:0] north5_out50;
wire [DATAWID-1:0] south5_out50;
wire [DATAWID-1:0] east5_out51;
wire [DATAWID-1:0] west5_out51;
wire [DATAWID-1:0] north5_out51;
wire [DATAWID-1:0] south5_out51;
wire [DATAWID-1:0] east5_out52;
wire [DATAWID-1:0] west5_out52;
wire [DATAWID-1:0] north5_out52;
wire [DATAWID-1:0] south5_out52;
wire [DATAWID-1:0] east5_out53;
wire [DATAWID-1:0] west5_out53;
wire [DATAWID-1:0] north5_out53;
wire [DATAWID-1:0] south5_out53;
wire [DATAWID-1:0] east5_out54;
wire [DATAWID-1:0] west5_out54;
wire [DATAWID-1:0] north5_out54;
wire [DATAWID-1:0] south5_out54;
wire [DATAWID-1:0] east5_out55;
wire [DATAWID-1:0] west5_out55;
wire [DATAWID-1:0] north5_out55;
wire [DATAWID-1:0] south5_out55;
wire [DATAWID-1:0] east5_out56;
wire [DATAWID-1:0] west5_out56;
wire [DATAWID-1:0] north5_out56;
wire [DATAWID-1:0] south5_out56;
wire [DATAWID-1:0] east5_out57;
wire [DATAWID-1:0] west5_out57;
wire [DATAWID-1:0] north5_out57;
wire [DATAWID-1:0] south5_out57;
wire [DATAWID-1:0] east5_out58;
wire [DATAWID-1:0] west5_out58;
wire [DATAWID-1:0] north5_out58;
wire [DATAWID-1:0] south5_out58;
wire [DATAWID-1:0] east5_out59;
wire [DATAWID-1:0] west5_out59;
wire [DATAWID-1:0] north5_out59;
wire [DATAWID-1:0] south5_out59;
wire [DATAWID-1:0] east6_out60;
wire [DATAWID-1:0] west6_out60;
wire [DATAWID-1:0] north6_out60;
wire [DATAWID-1:0] south6_out60;
wire [DATAWID-1:0] east6_out61;
wire [DATAWID-1:0] west6_out61;
wire [DATAWID-1:0] north6_out61;
wire [DATAWID-1:0] south6_out61;
wire [DATAWID-1:0] east6_out62;
wire [DATAWID-1:0] west6_out62;
wire [DATAWID-1:0] north6_out62;
wire [DATAWID-1:0] south6_out62;
wire [DATAWID-1:0] east6_out63;
wire [DATAWID-1:0] west6_out63;
wire [DATAWID-1:0] north6_out63;
wire [DATAWID-1:0] south6_out63;
wire [DATAWID-1:0] east6_out64;
wire [DATAWID-1:0] west6_out64;
wire [DATAWID-1:0] north6_out64;
wire [DATAWID-1:0] south6_out64;
wire [DATAWID-1:0] east6_out65;
wire [DATAWID-1:0] west6_out65;
wire [DATAWID-1:0] north6_out65;
wire [DATAWID-1:0] south6_out65;
wire [DATAWID-1:0] east6_out66;
wire [DATAWID-1:0] west6_out66;
wire [DATAWID-1:0] north6_out66;
wire [DATAWID-1:0] south6_out66;
wire [DATAWID-1:0] east6_out67;
wire [DATAWID-1:0] west6_out67;
wire [DATAWID-1:0] north6_out67;
wire [DATAWID-1:0] south6_out67;
wire [DATAWID-1:0] east6_out68;
wire [DATAWID-1:0] west6_out68;
wire [DATAWID-1:0] north6_out68;
wire [DATAWID-1:0] south6_out68;
wire [DATAWID-1:0] east6_out69;
wire [DATAWID-1:0] west6_out69;
wire [DATAWID-1:0] north6_out69;
wire [DATAWID-1:0] south6_out69;
wire [DATAWID-1:0] east7_out70;
wire [DATAWID-1:0] west7_out70;
wire [DATAWID-1:0] north7_out70;
wire [DATAWID-1:0] south7_out70;
wire [DATAWID-1:0] east7_out71;
wire [DATAWID-1:0] west7_out71;
wire [DATAWID-1:0] north7_out71;
wire [DATAWID-1:0] south7_out71;
wire [DATAWID-1:0] east7_out72;
wire [DATAWID-1:0] west7_out72;
wire [DATAWID-1:0] north7_out72;
wire [DATAWID-1:0] south7_out72;
wire [DATAWID-1:0] east7_out73;
wire [DATAWID-1:0] west7_out73;
wire [DATAWID-1:0] north7_out73;
wire [DATAWID-1:0] south7_out73;
wire [DATAWID-1:0] east7_out74;
wire [DATAWID-1:0] west7_out74;
wire [DATAWID-1:0] north7_out74;
wire [DATAWID-1:0] south7_out74;
wire [DATAWID-1:0] east7_out75;
wire [DATAWID-1:0] west7_out75;
wire [DATAWID-1:0] north7_out75;
wire [DATAWID-1:0] south7_out75;
wire [DATAWID-1:0] east7_out76;
wire [DATAWID-1:0] west7_out76;
wire [DATAWID-1:0] north7_out76;
wire [DATAWID-1:0] south7_out76;
wire [DATAWID-1:0] east7_out77;
wire [DATAWID-1:0] west7_out77;
wire [DATAWID-1:0] north7_out77;
wire [DATAWID-1:0] south7_out77;
wire [DATAWID-1:0] east7_out78;
wire [DATAWID-1:0] west7_out78;
wire [DATAWID-1:0] north7_out78;
wire [DATAWID-1:0] south7_out78;
wire [DATAWID-1:0] east7_out79;
wire [DATAWID-1:0] west7_out79;
wire [DATAWID-1:0] north7_out79;
wire [DATAWID-1:0] south7_out79;
wire [DATAWID-1:0] east8_out80;
wire [DATAWID-1:0] west8_out80;
wire [DATAWID-1:0] north8_out80;
wire [DATAWID-1:0] south8_out80;
wire [DATAWID-1:0] east8_out81;
wire [DATAWID-1:0] west8_out81;
wire [DATAWID-1:0] north8_out81;
wire [DATAWID-1:0] south8_out81;
wire [DATAWID-1:0] east8_out82;
wire [DATAWID-1:0] west8_out82;
wire [DATAWID-1:0] north8_out82;
wire [DATAWID-1:0] south8_out82;
wire [DATAWID-1:0] east8_out83;
wire [DATAWID-1:0] west8_out83;
wire [DATAWID-1:0] north8_out83;
wire [DATAWID-1:0] south8_out83;
wire [DATAWID-1:0] east8_out84;
wire [DATAWID-1:0] west8_out84;
wire [DATAWID-1:0] north8_out84;
wire [DATAWID-1:0] south8_out84;
wire [DATAWID-1:0] east8_out85;
wire [DATAWID-1:0] west8_out85;
wire [DATAWID-1:0] north8_out85;
wire [DATAWID-1:0] south8_out85;
wire [DATAWID-1:0] east8_out86;
wire [DATAWID-1:0] west8_out86;
wire [DATAWID-1:0] north8_out86;
wire [DATAWID-1:0] south8_out86;
wire [DATAWID-1:0] east8_out87;
wire [DATAWID-1:0] west8_out87;
wire [DATAWID-1:0] north8_out87;
wire [DATAWID-1:0] south8_out87;
wire [DATAWID-1:0] east8_out88;
wire [DATAWID-1:0] west8_out88;
wire [DATAWID-1:0] north8_out88;
wire [DATAWID-1:0] south8_out88;
wire [DATAWID-1:0] east8_out89;
wire [DATAWID-1:0] west8_out89;
wire [DATAWID-1:0] north8_out89;
wire [DATAWID-1:0] south8_out89;
wire [DATAWID-1:0] east9_out90;
wire [DATAWID-1:0] west9_out90;
wire [DATAWID-1:0] north9_out90;
wire [DATAWID-1:0] south9_out90;
wire [DATAWID-1:0] east9_out91;
wire [DATAWID-1:0] west9_out91;
wire [DATAWID-1:0] north9_out91;
wire [DATAWID-1:0] south9_out91;
wire [DATAWID-1:0] east9_out92;
wire [DATAWID-1:0] west9_out92;
wire [DATAWID-1:0] north9_out92;
wire [DATAWID-1:0] south9_out92;
wire [DATAWID-1:0] east9_out93;
wire [DATAWID-1:0] west9_out93;
wire [DATAWID-1:0] north9_out93;
wire [DATAWID-1:0] south9_out93;
wire [DATAWID-1:0] east9_out94;
wire [DATAWID-1:0] west9_out94;
wire [DATAWID-1:0] north9_out94;
wire [DATAWID-1:0] south9_out94;
wire [DATAWID-1:0] east9_out95;
wire [DATAWID-1:0] west9_out95;
wire [DATAWID-1:0] north9_out95;
wire [DATAWID-1:0] south9_out95;
wire [DATAWID-1:0] east9_out96;
wire [DATAWID-1:0] west9_out96;
wire [DATAWID-1:0] north9_out96;
wire [DATAWID-1:0] south9_out96;
wire [DATAWID-1:0] east9_out97;
wire [DATAWID-1:0] west9_out97;
wire [DATAWID-1:0] north9_out97;
wire [DATAWID-1:0] south9_out97;
wire [DATAWID-1:0] east9_out98;
wire [DATAWID-1:0] west9_out98;
wire [DATAWID-1:0] north9_out98;
wire [DATAWID-1:0] south9_out98;
wire [DATAWID-1:0] east9_out99;
wire [DATAWID-1:0] west9_out99;
wire [DATAWID-1:0] north9_out99;
wire [DATAWID-1:0] south9_out99;
router r000
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in00),
.i01(east0_in00),
.i02(west0_in00),
.i03(north0_in00),
.i04(south0_in00),
.o00(local0_out00),
.o01(east0_out00),
.o02(west0_out00),
.o03(north0_out00),
.o04(south0_out00)
);
router r001
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in01),
.i01(east0_in01),
.i02(west0_in01),
.i03(north0_in01),
.i04(south0_in01),
.o00(local0_out01),
.o01(east0_out01),
.o02(west0_out01),
.o03(north0_out01),
.o04(south0_out01)
);
router r002
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in02),
.i01(east0_in02),
.i02(west0_in02),
.i03(north0_in02),
.i04(south0_in02),
.o00(local0_out02),
.o01(east0_out02),
.o02(west0_out02),
.o03(north0_out02),
.o04(south0_out02)
);
router r003
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in03),
.i01(east0_in03),
.i02(west0_in03),
.i03(north0_in03),
.i04(south0_in03),
.o00(local0_out03),
.o01(east0_out03),
.o02(west0_out03),
.o03(north0_out03),
.o04(south0_out03)
);
router r004
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in04),
.i01(east0_in04),
.i02(west0_in04),
.i03(north0_in04),
.i04(south0_in04),
.o00(local0_out04),
.o01(east0_out04),
.o02(west0_out04),
.o03(north0_out04),
.o04(south0_out04)
);
router r005
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in05),
.i01(east0_in05),
.i02(west0_in05),
.i03(north0_in05),
.i04(south0_in05),
.o00(local0_out05),
.o01(east0_out05),
.o02(west0_out05),
.o03(north0_out05),
.o04(south0_out05)
);
router r006
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in06),
.i01(east0_in06),
.i02(west0_in06),
.i03(north0_in06),
.i04(south0_in06),
.o00(local0_out06),
.o01(east0_out06),
.o02(west0_out06),
.o03(north0_out06),
.o04(south0_out06)
);
router r007
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in07),
.i01(east0_in07),
.i02(west0_in07),
.i03(north0_in07),
.i04(south0_in07),
.o00(local0_out07),
.o01(east0_out07),
.o02(west0_out07),
.o03(north0_out07),
.o04(south0_out07)
);
router r008
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in08),
.i01(east0_in08),
.i02(west0_in08),
.i03(north0_in08),
.i04(south0_in08),
.o00(local0_out08),
.o01(east0_out08),
.o02(west0_out08),
.o03(north0_out08),
.o04(south0_out08)
);
router r009
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in09),
.i01(east0_in09),
.i02(west0_in09),
.i03(north0_in09),
.i04(south0_in09),
.o00(local0_out09),
.o01(east0_out09),
.o02(west0_out09),
.o03(north0_out09),
.o04(south0_out09)
);
router r110
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in10),
.i01(east1_in10),
.i02(west1_in10),
.i03(north1_in10),
.i04(south1_in10),
.o00(local1_out10),
.o01(east1_out10),
.o02(west1_out10),
.o03(north1_out10),
.o04(south1_out10)
);
router r111
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in11),
.i01(east1_in11),
.i02(west1_in11),
.i03(north1_in11),
.i04(south1_in11),
.o00(local1_out11),
.o01(east1_out11),
.o02(west1_out11),
.o03(north1_out11),
.o04(south1_out11)
);
router r112
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in12),
.i01(east1_in12),
.i02(west1_in12),
.i03(north1_in12),
.i04(south1_in12),
.o00(local1_out12),
.o01(east1_out12),
.o02(west1_out12),
.o03(north1_out12),
.o04(south1_out12)
);
router r113
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in13),
.i01(east1_in13),
.i02(west1_in13),
.i03(north1_in13),
.i04(south1_in13),
.o00(local1_out13),
.o01(east1_out13),
.o02(west1_out13),
.o03(north1_out13),
.o04(south1_out13)
);
router r114
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in14),
.i01(east1_in14),
.i02(west1_in14),
.i03(north1_in14),
.i04(south1_in14),
.o00(local1_out14),
.o01(east1_out14),
.o02(west1_out14),
.o03(north1_out14),
.o04(south1_out14)
);
router r115
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in15),
.i01(east1_in15),
.i02(west1_in15),
.i03(north1_in15),
.i04(south1_in15),
.o00(local1_out15),
.o01(east1_out15),
.o02(west1_out15),
.o03(north1_out15),
.o04(south1_out15)
);
router r116
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in16),
.i01(east1_in16),
.i02(west1_in16),
.i03(north1_in16),
.i04(south1_in16),
.o00(local1_out16),
.o01(east1_out16),
.o02(west1_out16),
.o03(north1_out16),
.o04(south1_out16)
);
router r117
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in17),
.i01(east1_in17),
.i02(west1_in17),
.i03(north1_in17),
.i04(south1_in17),
.o00(local1_out17),
.o01(east1_out17),
.o02(west1_out17),
.o03(north1_out17),
.o04(south1_out17)
);
router r118
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in18),
.i01(east1_in18),
.i02(west1_in18),
.i03(north1_in18),
.i04(south1_in18),
.o00(local1_out18),
.o01(east1_out18),
.o02(west1_out18),
.o03(north1_out18),
.o04(south1_out18)
);
router r119
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in19),
.i01(east1_in19),
.i02(west1_in19),
.i03(north1_in19),
.i04(south1_in19),
.o00(local1_out19),
.o01(east1_out19),
.o02(west1_out19),
.o03(north1_out19),
.o04(south1_out19)
);
router r220
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in20),
.i01(east2_in20),
.i02(west2_in20),
.i03(north2_in20),
.i04(south2_in20),
.o00(local2_out20),
.o01(east2_out20),
.o02(west2_out20),
.o03(north2_out20),
.o04(south2_out20)
);
router r221
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in21),
.i01(east2_in21),
.i02(west2_in21),
.i03(north2_in21),
.i04(south2_in21),
.o00(local2_out21),
.o01(east2_out21),
.o02(west2_out21),
.o03(north2_out21),
.o04(south2_out21)
);
router r222
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in22),
.i01(east2_in22),
.i02(west2_in22),
.i03(north2_in22),
.i04(south2_in22),
.o00(local2_out22),
.o01(east2_out22),
.o02(west2_out22),
.o03(north2_out22),
.o04(south2_out22)
);
router r223
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in23),
.i01(east2_in23),
.i02(west2_in23),
.i03(north2_in23),
.i04(south2_in23),
.o00(local2_out23),
.o01(east2_out23),
.o02(west2_out23),
.o03(north2_out23),
.o04(south2_out23)
);
router r224
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in24),
.i01(east2_in24),
.i02(west2_in24),
.i03(north2_in24),
.i04(south2_in24),
.o00(local2_out24),
.o01(east2_out24),
.o02(west2_out24),
.o03(north2_out24),
.o04(south2_out24)
);
router r225
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in25),
.i01(east2_in25),
.i02(west2_in25),
.i03(north2_in25),
.i04(south2_in25),
.o00(local2_out25),
.o01(east2_out25),
.o02(west2_out25),
.o03(north2_out25),
.o04(south2_out25)
);
router r226
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in26),
.i01(east2_in26),
.i02(west2_in26),
.i03(north2_in26),
.i04(south2_in26),
.o00(local2_out26),
.o01(east2_out26),
.o02(west2_out26),
.o03(north2_out26),
.o04(south2_out26)
);
router r227
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in27),
.i01(east2_in27),
.i02(west2_in27),
.i03(north2_in27),
.i04(south2_in27),
.o00(local2_out27),
.o01(east2_out27),
.o02(west2_out27),
.o03(north2_out27),
.o04(south2_out27)
);
router r228
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in28),
.i01(east2_in28),
.i02(west2_in28),
.i03(north2_in28),
.i04(south2_in28),
.o00(local2_out28),
.o01(east2_out28),
.o02(west2_out28),
.o03(north2_out28),
.o04(south2_out28)
);
router r229
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in29),
.i01(east2_in29),
.i02(west2_in29),
.i03(north2_in29),
.i04(south2_in29),
.o00(local2_out29),
.o01(east2_out29),
.o02(west2_out29),
.o03(north2_out29),
.o04(south2_out29)
);
router r330
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in30),
.i01(east3_in30),
.i02(west3_in30),
.i03(north3_in30),
.i04(south3_in30),
.o00(local3_out30),
.o01(east3_out30),
.o02(west3_out30),
.o03(north3_out30),
.o04(south3_out30)
);
router r331
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in31),
.i01(east3_in31),
.i02(west3_in31),
.i03(north3_in31),
.i04(south3_in31),
.o00(local3_out31),
.o01(east3_out31),
.o02(west3_out31),
.o03(north3_out31),
.o04(south3_out31)
);
router r332
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in32),
.i01(east3_in32),
.i02(west3_in32),
.i03(north3_in32),
.i04(south3_in32),
.o00(local3_out32),
.o01(east3_out32),
.o02(west3_out32),
.o03(north3_out32),
.o04(south3_out32)
);
router r333
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in33),
.i01(east3_in33),
.i02(west3_in33),
.i03(north3_in33),
.i04(south3_in33),
.o00(local3_out33),
.o01(east3_out33),
.o02(west3_out33),
.o03(north3_out33),
.o04(south3_out33)
);
router r334
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in34),
.i01(east3_in34),
.i02(west3_in34),
.i03(north3_in34),
.i04(south3_in34),
.o00(local3_out34),
.o01(east3_out34),
.o02(west3_out34),
.o03(north3_out34),
.o04(south3_out34)
);
router r335
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in35),
.i01(east3_in35),
.i02(west3_in35),
.i03(north3_in35),
.i04(south3_in35),
.o00(local3_out35),
.o01(east3_out35),
.o02(west3_out35),
.o03(north3_out35),
.o04(south3_out35)
);
router r336
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in36),
.i01(east3_in36),
.i02(west3_in36),
.i03(north3_in36),
.i04(south3_in36),
.o00(local3_out36),
.o01(east3_out36),
.o02(west3_out36),
.o03(north3_out36),
.o04(south3_out36)
);
router r337
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in37),
.i01(east3_in37),
.i02(west3_in37),
.i03(north3_in37),
.i04(south3_in37),
.o00(local3_out37),
.o01(east3_out37),
.o02(west3_out37),
.o03(north3_out37),
.o04(south3_out37)
);
router r338
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in38),
.i01(east3_in38),
.i02(west3_in38),
.i03(north3_in38),
.i04(south3_in38),
.o00(local3_out38),
.o01(east3_out38),
.o02(west3_out38),
.o03(north3_out38),
.o04(south3_out38)
);
router r339
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in39),
.i01(east3_in39),
.i02(west3_in39),
.i03(north3_in39),
.i04(south3_in39),
.o00(local3_out39),
.o01(east3_out39),
.o02(west3_out39),
.o03(north3_out39),
.o04(south3_out39)
);
router r440
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in40),
.i01(east4_in40),
.i02(west4_in40),
.i03(north4_in40),
.i04(south4_in40),
.o00(local4_out40),
.o01(east4_out40),
.o02(west4_out40),
.o03(north4_out40),
.o04(south4_out40)
);
router r441
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in41),
.i01(east4_in41),
.i02(west4_in41),
.i03(north4_in41),
.i04(south4_in41),
.o00(local4_out41),
.o01(east4_out41),
.o02(west4_out41),
.o03(north4_out41),
.o04(south4_out41)
);
router r442
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in42),
.i01(east4_in42),
.i02(west4_in42),
.i03(north4_in42),
.i04(south4_in42),
.o00(local4_out42),
.o01(east4_out42),
.o02(west4_out42),
.o03(north4_out42),
.o04(south4_out42)
);
router r443
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in43),
.i01(east4_in43),
.i02(west4_in43),
.i03(north4_in43),
.i04(south4_in43),
.o00(local4_out43),
.o01(east4_out43),
.o02(west4_out43),
.o03(north4_out43),
.o04(south4_out43)
);
router r444
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in44),
.i01(east4_in44),
.i02(west4_in44),
.i03(north4_in44),
.i04(south4_in44),
.o00(local4_out44),
.o01(east4_out44),
.o02(west4_out44),
.o03(north4_out44),
.o04(south4_out44)
);
router r445
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in45),
.i01(east4_in45),
.i02(west4_in45),
.i03(north4_in45),
.i04(south4_in45),
.o00(local4_out45),
.o01(east4_out45),
.o02(west4_out45),
.o03(north4_out45),
.o04(south4_out45)
);
router r446
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in46),
.i01(east4_in46),
.i02(west4_in46),
.i03(north4_in46),
.i04(south4_in46),
.o00(local4_out46),
.o01(east4_out46),
.o02(west4_out46),
.o03(north4_out46),
.o04(south4_out46)
);
router r447
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in47),
.i01(east4_in47),
.i02(west4_in47),
.i03(north4_in47),
.i04(south4_in47),
.o00(local4_out47),
.o01(east4_out47),
.o02(west4_out47),
.o03(north4_out47),
.o04(south4_out47)
);
router r448
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in48),
.i01(east4_in48),
.i02(west4_in48),
.i03(north4_in48),
.i04(south4_in48),
.o00(local4_out48),
.o01(east4_out48),
.o02(west4_out48),
.o03(north4_out48),
.o04(south4_out48)
);
router r449
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in49),
.i01(east4_in49),
.i02(west4_in49),
.i03(north4_in49),
.i04(south4_in49),
.o00(local4_out49),
.o01(east4_out49),
.o02(west4_out49),
.o03(north4_out49),
.o04(south4_out49)
);
router r550
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in50),
.i01(east5_in50),
.i02(west5_in50),
.i03(north5_in50),
.i04(south5_in50),
.o00(local5_out50),
.o01(east5_out50),
.o02(west5_out50),
.o03(north5_out50),
.o04(south5_out50)
);
router r551
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in51),
.i01(east5_in51),
.i02(west5_in51),
.i03(north5_in51),
.i04(south5_in51),
.o00(local5_out51),
.o01(east5_out51),
.o02(west5_out51),
.o03(north5_out51),
.o04(south5_out51)
);
router r552
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in52),
.i01(east5_in52),
.i02(west5_in52),
.i03(north5_in52),
.i04(south5_in52),
.o00(local5_out52),
.o01(east5_out52),
.o02(west5_out52),
.o03(north5_out52),
.o04(south5_out52)
);
router r553
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in53),
.i01(east5_in53),
.i02(west5_in53),
.i03(north5_in53),
.i04(south5_in53),
.o00(local5_out53),
.o01(east5_out53),
.o02(west5_out53),
.o03(north5_out53),
.o04(south5_out53)
);
router r554
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in54),
.i01(east5_in54),
.i02(west5_in54),
.i03(north5_in54),
.i04(south5_in54),
.o00(local5_out54),
.o01(east5_out54),
.o02(west5_out54),
.o03(north5_out54),
.o04(south5_out54)
);
router r555
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in55),
.i01(east5_in55),
.i02(west5_in55),
.i03(north5_in55),
.i04(south5_in55),
.o00(local5_out55),
.o01(east5_out55),
.o02(west5_out55),
.o03(north5_out55),
.o04(south5_out55)
);
router r556
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in56),
.i01(east5_in56),
.i02(west5_in56),
.i03(north5_in56),
.i04(south5_in56),
.o00(local5_out56),
.o01(east5_out56),
.o02(west5_out56),
.o03(north5_out56),
.o04(south5_out56)
);
router r557
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in57),
.i01(east5_in57),
.i02(west5_in57),
.i03(north5_in57),
.i04(south5_in57),
.o00(local5_out57),
.o01(east5_out57),
.o02(west5_out57),
.o03(north5_out57),
.o04(south5_out57)
);
router r558
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in58),
.i01(east5_in58),
.i02(west5_in58),
.i03(north5_in58),
.i04(south5_in58),
.o00(local5_out58),
.o01(east5_out58),
.o02(west5_out58),
.o03(north5_out58),
.o04(south5_out58)
);
router r559
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in59),
.i01(east5_in59),
.i02(west5_in59),
.i03(north5_in59),
.i04(south5_in59),
.o00(local5_out59),
.o01(east5_out59),
.o02(west5_out59),
.o03(north5_out59),
.o04(south5_out59)
);
router r660
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in60),
.i01(east6_in60),
.i02(west6_in60),
.i03(north6_in60),
.i04(south6_in60),
.o00(local6_out60),
.o01(east6_out60),
.o02(west6_out60),
.o03(north6_out60),
.o04(south6_out60)
);
router r661
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in61),
.i01(east6_in61),
.i02(west6_in61),
.i03(north6_in61),
.i04(south6_in61),
.o00(local6_out61),
.o01(east6_out61),
.o02(west6_out61),
.o03(north6_out61),
.o04(south6_out61)
);
router r662
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in62),
.i01(east6_in62),
.i02(west6_in62),
.i03(north6_in62),
.i04(south6_in62),
.o00(local6_out62),
.o01(east6_out62),
.o02(west6_out62),
.o03(north6_out62),
.o04(south6_out62)
);
router r663
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in63),
.i01(east6_in63),
.i02(west6_in63),
.i03(north6_in63),
.i04(south6_in63),
.o00(local6_out63),
.o01(east6_out63),
.o02(west6_out63),
.o03(north6_out63),
.o04(south6_out63)
);
router r664
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in64),
.i01(east6_in64),
.i02(west6_in64),
.i03(north6_in64),
.i04(south6_in64),
.o00(local6_out64),
.o01(east6_out64),
.o02(west6_out64),
.o03(north6_out64),
.o04(south6_out64)
);
router r665
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in65),
.i01(east6_in65),
.i02(west6_in65),
.i03(north6_in65),
.i04(south6_in65),
.o00(local6_out65),
.o01(east6_out65),
.o02(west6_out65),
.o03(north6_out65),
.o04(south6_out65)
);
router r666
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in66),
.i01(east6_in66),
.i02(west6_in66),
.i03(north6_in66),
.i04(south6_in66),
.o00(local6_out66),
.o01(east6_out66),
.o02(west6_out66),
.o03(north6_out66),
.o04(south6_out66)
);
router r667
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in67),
.i01(east6_in67),
.i02(west6_in67),
.i03(north6_in67),
.i04(south6_in67),
.o00(local6_out67),
.o01(east6_out67),
.o02(west6_out67),
.o03(north6_out67),
.o04(south6_out67)
);
router r668
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in68),
.i01(east6_in68),
.i02(west6_in68),
.i03(north6_in68),
.i04(south6_in68),
.o00(local6_out68),
.o01(east6_out68),
.o02(west6_out68),
.o03(north6_out68),
.o04(south6_out68)
);
router r669
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in69),
.i01(east6_in69),
.i02(west6_in69),
.i03(north6_in69),
.i04(south6_in69),
.o00(local6_out69),
.o01(east6_out69),
.o02(west6_out69),
.o03(north6_out69),
.o04(south6_out69)
);
router r770
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in70),
.i01(east7_in70),
.i02(west7_in70),
.i03(north7_in70),
.i04(south7_in70),
.o00(local7_out70),
.o01(east7_out70),
.o02(west7_out70),
.o03(north7_out70),
.o04(south7_out70)
);
router r771
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in71),
.i01(east7_in71),
.i02(west7_in71),
.i03(north7_in71),
.i04(south7_in71),
.o00(local7_out71),
.o01(east7_out71),
.o02(west7_out71),
.o03(north7_out71),
.o04(south7_out71)
);
router r772
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in72),
.i01(east7_in72),
.i02(west7_in72),
.i03(north7_in72),
.i04(south7_in72),
.o00(local7_out72),
.o01(east7_out72),
.o02(west7_out72),
.o03(north7_out72),
.o04(south7_out72)
);
router r773
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in73),
.i01(east7_in73),
.i02(west7_in73),
.i03(north7_in73),
.i04(south7_in73),
.o00(local7_out73),
.o01(east7_out73),
.o02(west7_out73),
.o03(north7_out73),
.o04(south7_out73)
);
router r774
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in74),
.i01(east7_in74),
.i02(west7_in74),
.i03(north7_in74),
.i04(south7_in74),
.o00(local7_out74),
.o01(east7_out74),
.o02(west7_out74),
.o03(north7_out74),
.o04(south7_out74)
);
router r775
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in75),
.i01(east7_in75),
.i02(west7_in75),
.i03(north7_in75),
.i04(south7_in75),
.o00(local7_out75),
.o01(east7_out75),
.o02(west7_out75),
.o03(north7_out75),
.o04(south7_out75)
);
router r776
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in76),
.i01(east7_in76),
.i02(west7_in76),
.i03(north7_in76),
.i04(south7_in76),
.o00(local7_out76),
.o01(east7_out76),
.o02(west7_out76),
.o03(north7_out76),
.o04(south7_out76)
);
router r777
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in77),
.i01(east7_in77),
.i02(west7_in77),
.i03(north7_in77),
.i04(south7_in77),
.o00(local7_out77),
.o01(east7_out77),
.o02(west7_out77),
.o03(north7_out77),
.o04(south7_out77)
);
router r778
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in78),
.i01(east7_in78),
.i02(west7_in78),
.i03(north7_in78),
.i04(south7_in78),
.o00(local7_out78),
.o01(east7_out78),
.o02(west7_out78),
.o03(north7_out78),
.o04(south7_out78)
);
router r779
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in79),
.i01(east7_in79),
.i02(west7_in79),
.i03(north7_in79),
.i04(south7_in79),
.o00(local7_out79),
.o01(east7_out79),
.o02(west7_out79),
.o03(north7_out79),
.o04(south7_out79)
);
router r880
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in80),
.i01(east8_in80),
.i02(west8_in80),
.i03(north8_in80),
.i04(south8_in80),
.o00(local8_out80),
.o01(east8_out80),
.o02(west8_out80),
.o03(north8_out80),
.o04(south8_out80)
);
router r881
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in81),
.i01(east8_in81),
.i02(west8_in81),
.i03(north8_in81),
.i04(south8_in81),
.o00(local8_out81),
.o01(east8_out81),
.o02(west8_out81),
.o03(north8_out81),
.o04(south8_out81)
);
router r882
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in82),
.i01(east8_in82),
.i02(west8_in82),
.i03(north8_in82),
.i04(south8_in82),
.o00(local8_out82),
.o01(east8_out82),
.o02(west8_out82),
.o03(north8_out82),
.o04(south8_out82)
);
router r883
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in83),
.i01(east8_in83),
.i02(west8_in83),
.i03(north8_in83),
.i04(south8_in83),
.o00(local8_out83),
.o01(east8_out83),
.o02(west8_out83),
.o03(north8_out83),
.o04(south8_out83)
);
router r884
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in84),
.i01(east8_in84),
.i02(west8_in84),
.i03(north8_in84),
.i04(south8_in84),
.o00(local8_out84),
.o01(east8_out84),
.o02(west8_out84),
.o03(north8_out84),
.o04(south8_out84)
);
router r885
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in85),
.i01(east8_in85),
.i02(west8_in85),
.i03(north8_in85),
.i04(south8_in85),
.o00(local8_out85),
.o01(east8_out85),
.o02(west8_out85),
.o03(north8_out85),
.o04(south8_out85)
);
router r886
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in86),
.i01(east8_in86),
.i02(west8_in86),
.i03(north8_in86),
.i04(south8_in86),
.o00(local8_out86),
.o01(east8_out86),
.o02(west8_out86),
.o03(north8_out86),
.o04(south8_out86)
);
router r887
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in87),
.i01(east8_in87),
.i02(west8_in87),
.i03(north8_in87),
.i04(south8_in87),
.o00(local8_out87),
.o01(east8_out87),
.o02(west8_out87),
.o03(north8_out87),
.o04(south8_out87)
);
router r888
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in88),
.i01(east8_in88),
.i02(west8_in88),
.i03(north8_in88),
.i04(south8_in88),
.o00(local8_out88),
.o01(east8_out88),
.o02(west8_out88),
.o03(north8_out88),
.o04(south8_out88)
);
router r889
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in89),
.i01(east8_in89),
.i02(west8_in89),
.i03(north8_in89),
.i04(south8_in89),
.o00(local8_out89),
.o01(east8_out89),
.o02(west8_out89),
.o03(north8_out89),
.o04(south8_out89)
);
router r990
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in90),
.i01(east9_in90),
.i02(west9_in90),
.i03(north9_in90),
.i04(south9_in90),
.o00(local9_out90),
.o01(east9_out90),
.o02(west9_out90),
.o03(north9_out90),
.o04(south9_out90)
);
router r991
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in91),
.i01(east9_in91),
.i02(west9_in91),
.i03(north9_in91),
.i04(south9_in91),
.o00(local9_out91),
.o01(east9_out91),
.o02(west9_out91),
.o03(north9_out91),
.o04(south9_out91)
);
router r992
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in92),
.i01(east9_in92),
.i02(west9_in92),
.i03(north9_in92),
.i04(south9_in92),
.o00(local9_out92),
.o01(east9_out92),
.o02(west9_out92),
.o03(north9_out92),
.o04(south9_out92)
);
router r993
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in93),
.i01(east9_in93),
.i02(west9_in93),
.i03(north9_in93),
.i04(south9_in93),
.o00(local9_out93),
.o01(east9_out93),
.o02(west9_out93),
.o03(north9_out93),
.o04(south9_out93)
);
router r994
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in94),
.i01(east9_in94),
.i02(west9_in94),
.i03(north9_in94),
.i04(south9_in94),
.o00(local9_out94),
.o01(east9_out94),
.o02(west9_out94),
.o03(north9_out94),
.o04(south9_out94)
);
router r995
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in95),
.i01(east9_in95),
.i02(west9_in95),
.i03(north9_in95),
.i04(south9_in95),
.o00(local9_out95),
.o01(east9_out95),
.o02(west9_out95),
.o03(north9_out95),
.o04(south9_out95)
);
router r996
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in96),
.i01(east9_in96),
.i02(west9_in96),
.i03(north9_in96),
.i04(south9_in96),
.o00(local9_out96),
.o01(east9_out96),
.o02(west9_out96),
.o03(north9_out96),
.o04(south9_out96)
);
router r997
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in97),
.i01(east9_in97),
.i02(west9_in97),
.i03(north9_in97),
.i04(south9_in97),
.o00(local9_out97),
.o01(east9_out97),
.o02(west9_out97),
.o03(north9_out97),
.o04(south9_out97)
);
router r998
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in98),
.i01(east9_in98),
.i02(west9_in98),
.i03(north9_in98),
.i04(south9_in98),
.o00(local9_out98),
.o01(east9_out98),
.o02(west9_out98),
.o03(north9_out98),
.o04(south9_out98)
);
router r999
( .clk(clk), .rst(reset),
.Read(Read),.Write(Write),.i00(local_in99),
.i01(east9_in99),
.i02(west9_in99),
.i03(north9_in99),
.i04(south9_in99),
.o00(local9_out99),
.o01(east9_out99),
.o02(west9_out99),
.o03(north9_out99),
.o04(south9_out99)
);
always @ ( posedge clk)
begin
west0_in01<=east0_out00;
east0_in09<=west0_out00;
south9_in90<=north0_out00;
north1_in10<=south0_out00;
west0_in02<=east0_out01;
east0_in00<=west0_out01;
north1_in11<=south0_out01;
south9_in91<=north0_out01;
west0_in03<=east0_out02;
east0_in01<=west0_out02;
north1_in12<=south0_out02;
south9_in92<=north0_out02;
west0_in04<=east0_out03;
east0_in02<=west0_out03;
north1_in13<=south0_out03;
south9_in93<=north0_out03;
west0_in05<=east0_out04;
east0_in03<=west0_out04;
north1_in14<=south0_out04;
south9_in94<=north0_out04;
west0_in06<=east0_out05;
east0_in04<=west0_out05;
north1_in15<=south0_out05;
south9_in95<=north0_out05;
west0_in07<=east0_out06;
east0_in05<=west0_out06;
north1_in16<=south0_out06;
south9_in96<=north0_out06;
west0_in08<=east0_out07;
east0_in06<=west0_out07;
north1_in17<=south0_out07;
south9_in97<=north0_out07;
west0_in09<=east0_out08;
east0_in07<=west0_out08;
north1_in18<=south0_out08;
south9_in98<=north0_out08;
west0_in00<=east0_out09;
east0_in08<=west0_out09;
north1_in19<=south0_out09;
south9_in99<=north0_out09;
west1_in11<=east1_out10;
east1_in19<=west1_out10;
north2_in20<=south1_out10;
south0_in00<=north1_out10;
west1_in12<=east1_out11;
east1_in10<=west1_out11;
south0_in01<=north1_out11;
north2_in21<=south1_out11;
west1_in13<=east1_out12;
east1_in11<=west1_out12;
south0_in02<=north1_out12;
north2_in22<=south1_out12;
west1_in14<=east1_out13;
east1_in12<=west1_out13;
south0_in03<=north1_out13;
north2_in23<=south1_out13;
west1_in15<=east1_out14;
east1_in13<=west1_out14;
south0_in04<=north1_out14;
north2_in24<=south1_out14;
west1_in16<=east1_out15;
east1_in14<=west1_out15;
south0_in05<=north1_out15;
north2_in25<=south1_out15;
west1_in17<=east1_out16;
east1_in15<=west1_out16;
south0_in06<=north1_out16;
north2_in26<=south1_out16;
west1_in18<=east1_out17;
east1_in16<=west1_out17;
south0_in07<=north1_out17;
north2_in27<=south1_out17;
west1_in19<=east1_out18;
east1_in17<=west1_out18;
south0_in08<=north1_out18;
north2_in28<=south1_out18;
west1_in10<=east1_out19;
east1_in18<=west1_out19;
north2_in29<=south1_out19;
south0_in09<=north1_out19;
west2_in21<=east2_out20;
east2_in29<=west2_out20;
north3_in30<=south2_out20;
south1_in10<=north2_out20;
west2_in22<=east2_out21;
east2_in20<=west2_out21;
south1_in11<=north2_out21;
north3_in31<=south2_out21;
west2_in23<=east2_out22;
east2_in21<=west2_out22;
south1_in12<=north2_out22;
north3_in32<=south2_out22;
west2_in24<=east2_out23;
east2_in22<=west2_out23;
south1_in13<=north2_out23;
north3_in33<=south2_out23;
west2_in25<=east2_out24;
east2_in23<=west2_out24;
south1_in14<=north2_out24;
north3_in34<=south2_out24;
west2_in26<=east2_out25;
east2_in24<=west2_out25;
south1_in15<=north2_out25;
north3_in35<=south2_out25;
west2_in27<=east2_out26;
east2_in25<=west2_out26;
south1_in16<=north2_out26;
north3_in36<=south2_out26;
west2_in28<=east2_out27;
east2_in26<=west2_out27;
south1_in17<=north2_out27;
north3_in37<=south2_out27;
west2_in29<=east2_out28;
east2_in27<=west2_out28;
south1_in18<=north2_out28;
north3_in38<=south2_out28;
west2_in20<=east2_out29;
east2_in28<=west2_out29;
north3_in39<=south2_out29;
south1_in19<=north2_out29;
west3_in31<=east3_out30;
east3_in39<=west3_out30;
north4_in40<=south3_out30;
south2_in20<=north3_out30;
west3_in32<=east3_out31;
east3_in30<=west3_out31;
south2_in21<=north3_out31;
north4_in41<=south3_out31;
west3_in33<=east3_out32;
east3_in31<=west3_out32;
south2_in22<=north3_out32;
north4_in42<=south3_out32;
west3_in34<=east3_out33;
east3_in32<=west3_out33;
south2_in23<=north3_out33;
north4_in43<=south3_out33;
west3_in35<=east3_out34;
east3_in33<=west3_out34;
south2_in24<=north3_out34;
north4_in44<=south3_out34;
west3_in36<=east3_out35;
east3_in34<=west3_out35;
south2_in25<=north3_out35;
north4_in45<=south3_out35;
west3_in37<=east3_out36;
east3_in35<=west3_out36;
south2_in26<=north3_out36;
north4_in46<=south3_out36;
west3_in38<=east3_out37;
east3_in36<=west3_out37;
south2_in27<=north3_out37;
north4_in47<=south3_out37;
west3_in39<=east3_out38;
east3_in37<=west3_out38;
south2_in28<=north3_out38;
north4_in48<=south3_out38;
west3_in30<=east3_out39;
east3_in38<=west3_out39;
north4_in49<=south3_out39;
south2_in29<=north3_out39;
west4_in41<=east4_out40;
east4_in49<=west4_out40;
north5_in50<=south4_out40;
south3_in30<=north4_out40;
west4_in42<=east4_out41;
east4_in40<=west4_out41;
south3_in31<=north4_out41;
north5_in51<=south4_out41;
west4_in43<=east4_out42;
east4_in41<=west4_out42;
south3_in32<=north4_out42;
north5_in52<=south4_out42;
west4_in44<=east4_out43;
east4_in42<=west4_out43;
south3_in33<=north4_out43;
north5_in53<=south4_out43;
west4_in45<=east4_out44;
east4_in43<=west4_out44;
south3_in34<=north4_out44;
north5_in54<=south4_out44;
west4_in46<=east4_out45;
east4_in44<=west4_out45;
south3_in35<=north4_out45;
north5_in55<=south4_out45;
west4_in47<=east4_out46;
east4_in45<=west4_out46;
south3_in36<=north4_out46;
north5_in56<=south4_out46;
west4_in48<=east4_out47;
east4_in46<=west4_out47;
south3_in37<=north4_out47;
north5_in57<=south4_out47;
west4_in49<=east4_out48;
east4_in47<=west4_out48;
south3_in38<=north4_out48;
north5_in58<=south4_out48;
west4_in40<=east4_out49;
east4_in48<=west4_out49;
north5_in59<=south4_out49;
south3_in39<=north4_out49;
west5_in51<=east5_out50;
east5_in59<=west5_out50;
north6_in60<=south5_out50;
south4_in40<=north5_out50;
west5_in52<=east5_out51;
east5_in50<=west5_out51;
south4_in41<=north5_out51;
north6_in61<=south5_out51;
west5_in53<=east5_out52;
east5_in51<=west5_out52;
south4_in42<=north5_out52;
north6_in62<=south5_out52;
west5_in54<=east5_out53;
east5_in52<=west5_out53;
south4_in43<=north5_out53;
north6_in63<=south5_out53;
west5_in55<=east5_out54;
east5_in53<=west5_out54;
south4_in44<=north5_out54;
north6_in64<=south5_out54;
west5_in56<=east5_out55;
east5_in54<=west5_out55;
south4_in45<=north5_out55;
north6_in65<=south5_out55;
west5_in57<=east5_out56;
east5_in55<=west5_out56;
south4_in46<=north5_out56;
north6_in66<=south5_out56;
west5_in58<=east5_out57;
east5_in56<=west5_out57;
south4_in47<=north5_out57;
north6_in67<=south5_out57;
west5_in59<=east5_out58;
east5_in57<=west5_out58;
south4_in48<=north5_out58;
north6_in68<=south5_out58;
west5_in50<=east5_out59;
east5_in58<=west5_out59;
north6_in69<=south5_out59;
south4_in49<=north5_out59;
west6_in61<=east6_out60;
east6_in69<=west6_out60;
north7_in70<=south6_out60;
south5_in50<=north6_out60;
west6_in62<=east6_out61;
east6_in60<=west6_out61;
south5_in51<=north6_out61;
north7_in71<=south6_out61;
west6_in63<=east6_out62;
east6_in61<=west6_out62;
south5_in52<=north6_out62;
north7_in72<=south6_out62;
west6_in64<=east6_out63;
east6_in62<=west6_out63;
south5_in53<=north6_out63;
north7_in73<=south6_out63;
west6_in65<=east6_out64;
east6_in63<=west6_out64;
south5_in54<=north6_out64;
north7_in74<=south6_out64;
west6_in66<=east6_out65;
east6_in64<=west6_out65;
south5_in55<=north6_out65;
north7_in75<=south6_out65;
west6_in67<=east6_out66;
east6_in65<=west6_out66;
south5_in56<=north6_out66;
north7_in76<=south6_out66;
west6_in68<=east6_out67;
east6_in66<=west6_out67;
south5_in57<=north6_out67;
north7_in77<=south6_out67;
west6_in69<=east6_out68;
east6_in67<=west6_out68;
south5_in58<=north6_out68;
north7_in78<=south6_out68;
west6_in60<=east6_out69;
east6_in68<=west6_out69;
north7_in79<=south6_out69;
south5_in59<=north6_out69;
west7_in71<=east7_out70;
east7_in79<=west7_out70;
north8_in80<=south7_out70;
south6_in60<=north7_out70;
west7_in72<=east7_out71;
east7_in70<=west7_out71;
south6_in61<=north7_out71;
north8_in81<=south7_out71;
west7_in73<=east7_out72;
east7_in71<=west7_out72;
south6_in62<=north7_out72;
north8_in82<=south7_out72;
west7_in74<=east7_out73;
east7_in72<=west7_out73;
south6_in63<=north7_out73;
north8_in83<=south7_out73;
west7_in75<=east7_out74;
east7_in73<=west7_out74;
south6_in64<=north7_out74;
north8_in84<=south7_out74;
west7_in76<=east7_out75;
east7_in74<=west7_out75;
south6_in65<=north7_out75;
north8_in85<=south7_out75;
west7_in77<=east7_out76;
east7_in75<=west7_out76;
south6_in66<=north7_out76;
north8_in86<=south7_out76;
west7_in78<=east7_out77;
east7_in76<=west7_out77;
south6_in67<=north7_out77;
north8_in87<=south7_out77;
west7_in79<=east7_out78;
east7_in77<=west7_out78;
south6_in68<=north7_out78;
north8_in88<=south7_out78;
west7_in70<=east7_out79;
east7_in78<=west7_out79;
north8_in89<=south7_out79;
south6_in69<=north7_out79;
west8_in81<=east8_out80;
east8_in89<=west8_out80;
north9_in90<=south8_out80;
south7_in70<=north8_out80;
west8_in82<=east8_out81;
east8_in80<=west8_out81;
south7_in71<=north8_out81;
north9_in91<=south8_out81;
west8_in83<=east8_out82;
east8_in81<=west8_out82;
south7_in72<=north8_out82;
north9_in92<=south8_out82;
west8_in84<=east8_out83;
east8_in82<=west8_out83;
south7_in73<=north8_out83;
north9_in93<=south8_out83;
west8_in85<=east8_out84;
east8_in83<=west8_out84;
south7_in74<=north8_out84;
north9_in94<=south8_out84;
west8_in86<=east8_out85;
east8_in84<=west8_out85;
south7_in75<=north8_out85;
north9_in95<=south8_out85;
west8_in87<=east8_out86;
east8_in85<=west8_out86;
south7_in76<=north8_out86;
north9_in96<=south8_out86;
west8_in88<=east8_out87;
east8_in86<=west8_out87;
south7_in77<=north8_out87;
north9_in97<=south8_out87;
west8_in89<=east8_out88;
east8_in87<=west8_out88;
south7_in78<=north8_out88;
north9_in98<=south8_out88;
west8_in80<=east8_out89;
east8_in88<=west8_out89;
north9_in99<=south8_out89;
south7_in79<=north8_out89;
west9_in91<=east9_out90;
east9_in99<=west9_out90;
north0_in00<=south9_out90;
south8_in80<=north9_out90;
west9_in92<=east9_out91;
east9_in90<=west9_out91;
south0_in01<=south9_out91;
south8_in81<=north9_out91;
west9_in93<=east9_out92;
east9_in91<=west9_out92;
south0_in02<=south9_out92;
south8_in82<=north9_out92;
west9_in94<=east9_out93;
east9_in92<=west9_out93;
south0_in03<=south9_out93;
south8_in83<=north9_out93;
west9_in95<=east9_out94;
east9_in93<=west9_out94;
south0_in04<=south9_out94;
south8_in84<=north9_out94;
west9_in96<=east9_out95;
east9_in94<=west9_out95;
south0_in05<=south9_out95;
south8_in85<=north9_out95;
west9_in97<=east9_out96;
east9_in95<=west9_out96;
south0_in06<=south9_out96;
south8_in86<=north9_out96;
west9_in98<=east9_out97;
east9_in96<=west9_out97;
south0_in07<=south9_out97;
south8_in87<=north9_out97;
west9_in99<=east9_out98;
east9_in97<=west9_out98;
south0_in08<=south9_out98;
south8_in88<=north9_out98;
west9_in90<=east9_out99;
east9_in98<=west9_out99;
north0_in09<=south9_out99;
south8_in89<=north9_out99;
end
endmodule
