`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    18:15:35 08/25/2016 
// Design Name: 
// Module Name:    crossbar 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module crossbar(i0,i1,i2,i3,i4,i5,i6,i7,i8,i9, i10, i11,i12,i13, i14,
      sel0, sel1,sel2,sel3,sel4, sel5,sel6,sel7,sel8,sel9,sel10, sel11,sel12,sel13,sel14,
      o0,o1,o2,o3,o4,o5,o6,o7,o8,o9,o10, o11,o12,o13,o14, clk, rst
    );
input clk, rst;
input[7:0] i0,i1,i2,i3,i4,i5,i6,i7,i8,i9, i10, i11,i12,i13, i14;
output reg[7:0] oo0,o1,o2,o3,o4,o5,o6,o7,o8,o9,o10, o11,o12,o13,o14;
input[9:0] sel0, sel1,sel2,sel3,sel4, sel5,sel6,sel7,sel8,sel9,sel10, sel11,sel12,sel13,sel14;
always @(posedge clk)
begin
case(sel0)
15'b000000000000001: o0<=i0;
15'b000000000000010: o0<=i1;
15'b000000000000100: o0<=i2;
15'b000000000001000: o0<=i3;
15'b000000000010000: o0<=i4;
15'b000000000100000: o0<=i5;
15'b000000001000000: o0<=i6;
15'b000000010000000: o0<=i7;
15'b000000100000000: o0<=i8;
15'b000001000000000: o0<=i9;
15'b000010000000000: o0<=i10;
15'b000100000000000: o0<=i11;
15'b001000000000000: o0<=i12;
15'b010000000000000: o0<=i13;
15'b100000000000000: o0<=i14;
default: o0<=15'bxxxxxxxxxxxxx;
endcase
case(sel1)
15'b000000000000001: o1<=i0;
15'b000000000000010: o1<=i1;
15'b000000000000100: o1<=i2;
15'b000000000001000: o1<=i3;
15'b000000000010000: o1<=i4;
15'b000000000100000: o1<=i5;
15'b000000001000000: o1<=i6;
15'b000000010000000: o1<=i7;
15'b000000100000000: o1<=i8;
15'b000001000000000: o1<=i9;
15'b000010000000000: o1<=i10;
15'b000100000000000: o1<=i11;
15'b001000000000000: o1<=i12;
15'b010000000000000: o1<=i13;
15'b100000000000000: o1<=i14;
default: o1<=15'bxxxxxxxxxxxxx;
endcase
case(sel2)
15'b000000000000001: o2<=i0;
15'b000000000000010: o2<=i1;
15'b000000000000100: o2<=i2;
15'b000000000001000: o2<=i3;
15'b000000000010000: o2<=i4;
15'b000000000100000: o2<=i5;
15'b000000001000000: o2<=i6;
15'b000000010000000: o2<=i7;
15'b000000100000000: o2<=i8;
15'b000001000000000: o2<=i9;
15'b000010000000000: o2<=i10;
15'b000100000000000: o2<=i11;
15'b001000000000000: o2<=i12;
15'b010000000000000: o2<=i13;
15'b100000000000000: o2<=i14;
default: o2<=15'bxxxxxxxxxxxxx;
endcase
case(sel3)
15'b000000000000001: o3<=i0;
15'b000000000000010: o3<=i1;
15'b000000000000100: o3<=i2;
15'b000000000001000: o3<=i3;
15'b000000000010000: o3<=i4;
15'b000000000100000: o3<=i5;
15'b000000001000000: o3<=i6;
15'b000000010000000: o3<=i7;
15'b000000100000000: o3<=i8;
15'b000001000000000: o3<=i9;
15'b000010000000000: o3<=i10;
15'b000100000000000: o3<=i11;
15'b001000000000000: o3<=i12;
15'b010000000000000: o3<=i13;
15'b100000000000000: o3<=i14;
default: o3<=15'bxxxxxxxxxxxxx;
endcase
case(sel4)
15'b000000000000001: o4<=i0;
15'b000000000000010: o4<=i1;
15'b000000000000100: o4<=i2;
15'b000000000001000: o4<=i3;
15'b000000000010000: o4<=i4;
15'b000000000100000: o4<=i5;
15'b000000001000000: o4<=i6;
15'b000000010000000: o4<=i7;
15'b000000100000000: o4<=i8;
15'b000001000000000: o4<=i9;
15'b000010000000000: o4<=i10;
15'b000100000000000: o4<=i11;
15'b001000000000000: o4<=i12;
15'b010000000000000: o4<=i13;
15'b100000000000000: o4<=i14;
default: o4<=15'bxxxxxxxxxxxxx;
endcase
case(sel5)
15'b000000000000001: o5<=i0;
15'b000000000000010: o5<=i1;
15'b000000000000100: o5<=i2;
15'b000000000001000: o5<=i3;
15'b000000000010000: o5<=i4;
15'b000000000100000: o5<=i5;
15'b000000001000000: o5<=i6;
15'b000000010000000: o5<=i7;
15'b000000100000000: o5<=i8;
15'b000001000000000: o5<=i9;
15'b000010000000000: o5<=i10;
15'b000100000000000: o5<=i11;
15'b001000000000000: o5<=i12;
15'b010000000000000: o5<=i13;
15'b100000000000000: o5<=i14;
default: o5<=15'bxxxxxxxxxxxxx;
endcase
case(sel6)
15'b000000000000001: o6<=i0;
15'b000000000000010: o6<=i1;
15'b000000000000100: o6<=i2;
15'b000000000001000: o6<=i3;
15'b000000000010000: o6<=i4;
15'b000000000100000: o6<=i5;
15'b000000001000000: o6<=i6;
15'b000000010000000: o6<=i7;
15'b000000100000000: o6<=i8;
15'b000001000000000: o6<=i9;
15'b000010000000000: o6<=i10;
15'b000100000000000: o6<=i11;
15'b001000000000000: o6<=i12;
15'b010000000000000: o6<=i13;
15'b100000000000000: o6<=i14;
default: o6<=15'bxxxxxxxxxxxxx;
endcase
case(sel7)
15'b000000000000001: o7<=i0;
15'b000000000000010: o7<=i1;
15'b000000000000100: o7<=i2;
15'b000000000001000: o7<=i3;
15'b000000000010000: o7<=i4;
15'b000000000100000: o7<=i5;
15'b000000001000000: o7<=i6;
15'b000000010000000: o7<=i7;
15'b000000100000000: o7<=i8;
15'b000001000000000: o7<=i9;
15'b000010000000000: o7<=i10;
15'b000100000000000: o7<=i11;
15'b001000000000000: o7<=i12;
15'b010000000000000: o7<=i13;
15'b100000000000000: o7<=i14;
default: o7<=15'bxxxxxxxxxxxxx;
endcase
case(sel8)
15'b000000000000001: o8<=i0;
15'b000000000000010: o8<=i1;
15'b000000000000100: o8<=i2;
15'b000000000001000: o8<=i3;
15'b000000000010000: o8<=i4;
15'b000000000100000: o8<=i5;
15'b000000001000000: o8<=i6;
15'b000000010000000: o8<=i7;
15'b000000100000000: o8<=i8;
15'b000001000000000: o8<=i9;
15'b000010000000000: o8<=i10;
15'b000100000000000: o8<=i11;
15'b001000000000000: o8<=i12;
15'b010000000000000: o8<=i13;
15'b100000000000000: o8<=i14;
default: o8<=15'bxxxxxxxxxxxxx;
endcase
case(sel9)
15'b000000000000001: o9<=i0;
15'b000000000000010: o9<=i1;
15'b000000000000100: o9<=i2;
15'b000000000001000: o9<=i3;
15'b000000000010000: o9<=i4;
15'b000000000100000: o9<=i5;
15'b000000001000000: o9<=i6;
15'b000000010000000: o9<=i7;
15'b000000100000000: o9<=i8;
15'b000001000000000: o9<=i9;
15'b000010000000000: o9<=i10;
15'b000100000000000: o9<=i11;
15'b001000000000000: o9<=i12;
15'b010000000000000: o9<=i13;
15'b100000000000000: o9<=i14;
default: o9<=15'bxxxxxxxxxxxxx;
endcase
case(sel10)
15'b000000000000001: o10<=i0;
15'b000000000000010: o10<=i1;
15'b000000000000100: o10<=i2;
15'b000000000001000: o10<=i3;
15'b000000000010000: o10<=i4;
15'b000000000100000: o10<=i5;
15'b000000001000000: o10<=i6;
15'b000000010000000: o10<=i7;
15'b000000100000000: o10<=i8;
15'b000001000000000: o10<=i9;
15'b000010000000000: o10<=i10;
15'b000100000000000: o10<=i11;
15'b001000000000000: o10<=i12;
15'b010000000000000: o10<=i13;
15'b100000000000000: o10<=i14;
default: o10<=15'bxxxxxxxxxxxxx;
endcase
case(sel11)
15'b000000000000001: o11<=i0;
15'b000000000000010: o11<=i1;
15'b000000000000100: o11<=i2;
15'b000000000001000: o11<=i3;
15'b000000000010000: o11<=i4;
15'b000000000100000: o11<=i5;
15'b000000001000000: o11<=i6;
15'b000000010000000: o11<=i7;
15'b000000100000000: o11<=i8;
15'b000001000000000: o11<=i9;
15'b000010000000000: o11<=i10;
15'b000100000000000: o11<=i11;
15'b001000000000000: o11<=i12;
15'b010000000000000: o11<=i13;
15'b100000000000000: o11<=i14;
default: o11<=15'bxxxxxxxxxxxxx;
endcase
case(sel12)
15'b000000000000001: o12<=i0;
15'b000000000000010: o12<=i1;
15'b000000000000100: o12<=i2;
15'b000000000001000: o12<=i3;
15'b000000000010000: o12<=i4;
15'b000000000100000: o12<=i5;
15'b000000001000000: o12<=i6;
15'b000000010000000: o12<=i7;
15'b000000100000000: o12<=i8;
15'b000001000000000: o12<=i9;
15'b000010000000000: o12<=i10;
15'b000100000000000: o12<=i11;
15'b001000000000000: o12<=i12;
15'b010000000000000: o12<=i13;
15'b100000000000000: o12<=i14;
default: o12<=15'bxxxxxxxxxxxxx;
endcase
case(sel13)
15'b000000000000001: o13<=i0;
15'b000000000000010: o13<=i1;
15'b000000000000100: o13<=i2;
15'b000000000001000: o13<=i3;
15'b000000000010000: o13<=i4;
15'b000000000100000: o13<=i5;
15'b000000001000000: o13<=i6;
15'b000000010000000: o13<=i7;
15'b000000100000000: o13<=i8;
15'b000001000000000: o13<=i9;
15'b000010000000000: o13<=i10;
15'b000100000000000: o13<=i11;
15'b001000000000000: o13<=i12;
15'b010000000000000: o13<=i13;
15'b100000000000000: o13<=i14;
default: o13<=15'bxxxxxxxxxxxxx;
endcase
case(sel14)
15'b000000000000001: o14<=i0;
15'b000000000000010: o14<=i1;
15'b000000000000100: o14<=i2;
15'b000000000001000: o14<=i3;
15'b000000000010000: o14<=i4;
15'b000000000100000: o14<=i5;
15'b000000001000000: o14<=i6;
15'b000000010000000: o14<=i7;
15'b000000100000000: o14<=i8;
15'b000001000000000: o14<=i9;
15'b000010000000000: o14<=i10;
15'b000100000000000: o14<=i11;
15'b001000000000000: o14<=i12;
15'b010000000000000: o14<=i13;
15'b100000000000000: o14<=i14;
default: o14<=15'bxxxxxxxxxxxxx;
endcase
$display("output local i0 %d, %t", i0, $time);
$display("output local i1 %d, %t", i1, $time);
$display("output local i2 %d, %t", i2, $time);
$display("output local i3 %d, %t", i3, $time);
$display("output local i4 %d, %t", i4, $time);
$display("select0 signal %b, %t", sel0, $time);
$display("select1 signal %b, %t", sel1, $time);
$display("select2 signal %b, %t", sel2, $time);
$display("select3 signal %b, %t", sel3, $time);
$display("select4 signal %b, %t", sel4, $time);


end
//sel1,sel2,sel3,sel4;
//assign o0= (i0&sel0);
//assign o0=((i0&~i1&~i2&~i3&~i4&sel0)|(~i0&i1&~i2&~i3&~i4&sel0)|(~i0&~i1&i2&~i3&~i4&sel0)|(~i0&~i1&~i2&i3&~i4&sel0)|(~i0&~i1&~i2&~i3&i4&sel0));
//assign o1=((i0&~i1&~i2&~i3&~i4&sel1)|(~i0&i1&~i2&~i3&~i4&sel1)|(~i0&~i1&i2&~i3&~i4&sel1)|(~i0&~i1&~i2&i3&~i4&sel1)|(~i0&~i1&~i2&~i3&i4&sel1));
//assign o2=((i0&~i1&~i2&~i3&~i4&sel2)|(~i0&i1&~i2&~i3&~i4&sel2)|(~i0&~i1&i2&~i3&~i4&sel2)|(~i0&~i1&~i2&i3&~i4&sel2)|(~i0&~i1&~i2&~i3&i4&sel2));
//assign o3=((i0&~i1&~i2&~i3&~i4&sel3)|(~i0&i1&~i2&~i3&~i4&sel3)|(~i0&~i1&i2&~i3&~i4&sel3)|(~i0&~i1&~i2&i3&~i4&sel3)|(~i0&~i1&~i2&~i3&i4&sel3));
//assign o4=((i0&~i1&~i2&~i3&~i4&sel4)|(~i0&i1&~i2&~i3&~i4&sel4)|(~i0&~i1&i2&~i3&~i4&sel4)|(~i0&~i1&~i2&i3&~i4&sel4)|(~i0&~i1&~i2&~i3&i4&sel4));
endmodule



