module test_case_0 #(parameter NUM_AGENT=6,
                     parameter PIPE_DLY =4,
                     parameter N = 10,
                     parameter M = 20
                    ) 
                    (
                         input  logic                 clk,
                         input  logic                 rst_n,
                         input  logic [NUM_AGENT-1:0] req,
                         output logic [NUM_AGENT-1:0] gnt,
                         output logic [2:0]           arbiter_state,
                         output logic                 arb_idle,
                         output logic                 arb_busy
                         abc.xyz [NUM_AGENT:0] arb_unbusy [1:8]
                    ) ;
bla bla
bla bla
bla bla
bla bla
bla bla
bla bla
bla bla
bla bla
bla bla
bla bla
endmodule
